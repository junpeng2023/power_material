module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net1028;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net1032;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net1033;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire clknet_0_clk;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net1021;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1029;
 wire net1030;
 wire net1031;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net914;
 wire clknet_1_0__leaf_net914;
 wire clknet_1_1__leaf_net914;
 wire clknet_0_net548;
 wire clknet_1_0__leaf_net548;
 wire clknet_1_1__leaf_net548;
 wire clknet_0_net666;
 wire clknet_1_0__leaf_net666;
 wire clknet_1_1__leaf_net666;
 wire clknet_0_net665;
 wire clknet_1_0__leaf_net665;
 wire clknet_1_1__leaf_net665;
 wire clknet_0_net894;
 wire clknet_1_0__leaf_net894;
 wire clknet_1_1__leaf_net894;
 wire clknet_0_net724;
 wire clknet_1_0__leaf_net724;
 wire clknet_1_1__leaf_net724;
 wire clknet_0_net715;
 wire clknet_1_0__leaf_net715;
 wire clknet_1_1__leaf_net715;
 wire clknet_0_net711;
 wire clknet_1_0__leaf_net711;
 wire clknet_1_1__leaf_net711;
 wire clknet_0_net655;
 wire clknet_1_0__leaf_net655;
 wire clknet_1_1__leaf_net655;
 wire clknet_0_net657;
 wire clknet_1_0__leaf_net657;
 wire clknet_1_1__leaf_net657;
 wire clknet_0_net912;
 wire clknet_1_0__leaf_net912;
 wire clknet_1_1__leaf_net912;
 wire clknet_0_net662;
 wire clknet_1_0__leaf_net662;
 wire clknet_1_1__leaf_net662;
 wire clknet_0_net664;
 wire clknet_1_0__leaf_net664;
 wire clknet_1_1__leaf_net664;
 wire clknet_0_net409;
 wire clknet_1_0__leaf_net409;
 wire clknet_1_1__leaf_net409;
 wire clknet_0_net460;
 wire clknet_1_0__leaf_net460;
 wire clknet_1_1__leaf_net460;
 wire clknet_0_net467;
 wire clknet_1_0__leaf_net467;
 wire clknet_1_1__leaf_net467;
 wire clknet_0_net466;
 wire clknet_1_0__leaf_net466;
 wire clknet_1_1__leaf_net466;
 wire clknet_0_net593;
 wire clknet_1_0__leaf_net593;
 wire clknet_1_1__leaf_net593;
 wire clknet_0_net583;
 wire clknet_1_0__leaf_net583;
 wire clknet_1_1__leaf_net583;
 wire clknet_0_net464;
 wire clknet_1_0__leaf_net464;
 wire clknet_1_1__leaf_net464;
 wire clknet_0_net728;
 wire clknet_1_0__leaf_net728;
 wire clknet_1_1__leaf_net728;
 wire clknet_0_net581;
 wire clknet_1_0__leaf_net581;
 wire clknet_1_1__leaf_net581;
 wire clknet_0_net957;
 wire clknet_1_0__leaf_net957;
 wire clknet_1_1__leaf_net957;
 wire clknet_0_net580;
 wire clknet_1_0__leaf_net580;
 wire clknet_1_1__leaf_net580;
 wire clknet_0_net472;
 wire clknet_1_0__leaf_net472;
 wire clknet_1_1__leaf_net472;
 wire clknet_0_net461;
 wire clknet_1_0__leaf_net461;
 wire clknet_1_1__leaf_net461;
 wire clknet_0_net621;
 wire clknet_1_0__leaf_net621;
 wire clknet_1_1__leaf_net621;
 wire clknet_0_net613;
 wire clknet_1_0__leaf_net613;
 wire clknet_1_1__leaf_net613;
 wire clknet_0_net611;
 wire clknet_1_0__leaf_net611;
 wire clknet_1_1__leaf_net611;
 wire clknet_0_net486;
 wire clknet_1_0__leaf_net486;
 wire clknet_1_1__leaf_net486;
 wire clknet_0_net459;
 wire clknet_1_0__leaf_net459;
 wire clknet_1_1__leaf_net459;
 wire clknet_0_net822;
 wire clknet_1_0__leaf_net822;
 wire clknet_1_1__leaf_net822;
 wire clknet_0_net427;
 wire clknet_1_0__leaf_net427;
 wire clknet_1_1__leaf_net427;
 wire clknet_0_net430;
 wire clknet_1_0__leaf_net430;
 wire clknet_1_1__leaf_net430;
 wire clknet_0_net420;
 wire clknet_1_0__leaf_net420;
 wire clknet_1_1__leaf_net420;
 wire clknet_0_net554;
 wire clknet_1_0__leaf_net554;
 wire clknet_1_1__leaf_net554;
 wire clknet_0_net678;
 wire clknet_1_0__leaf_net678;
 wire clknet_1_1__leaf_net678;
 wire clknet_0_net696;
 wire clknet_1_0__leaf_net696;
 wire clknet_1_1__leaf_net696;
 wire clknet_0_net557;
 wire clknet_1_0__leaf_net557;
 wire clknet_1_1__leaf_net557;
 wire clknet_0_net579;
 wire clknet_1_0__leaf_net579;
 wire clknet_1_1__leaf_net579;
 wire clknet_0_net913;
 wire clknet_1_0__leaf_net913;
 wire clknet_1_1__leaf_net913;
 wire clknet_0_net234;
 wire clknet_1_0__leaf_net234;
 wire clknet_1_1__leaf_net234;
 wire clknet_0_net240;
 wire clknet_1_0__leaf_net240;
 wire clknet_1_1__leaf_net240;
 wire clknet_0_net841;
 wire clknet_1_0__leaf_net841;
 wire clknet_1_1__leaf_net841;
 wire clknet_0_net499;
 wire clknet_1_0__leaf_net499;
 wire clknet_1_1__leaf_net499;
 wire clknet_0_net502;
 wire clknet_1_0__leaf_net502;
 wire clknet_1_1__leaf_net502;
 wire clknet_0_net875;
 wire clknet_1_0__leaf_net875;
 wire clknet_1_1__leaf_net875;
 wire clknet_0_net214;
 wire clknet_1_0__leaf_net214;
 wire clknet_1_1__leaf_net214;
 wire clknet_0_net858;
 wire clknet_1_0__leaf_net858;
 wire clknet_1_1__leaf_net858;
 wire clknet_0_net223;
 wire clknet_1_0__leaf_net223;
 wire clknet_1_1__leaf_net223;
 wire clknet_0_net241;
 wire clknet_1_0__leaf_net241;
 wire clknet_1_1__leaf_net241;
 wire clknet_0_net839;
 wire clknet_1_0__leaf_net839;
 wire clknet_1_1__leaf_net839;
 wire clknet_0_net222;
 wire clknet_1_0__leaf_net222;
 wire clknet_1_1__leaf_net222;
 wire clknet_0_net352;
 wire clknet_1_0__leaf_net352;
 wire clknet_1_1__leaf_net352;
 wire clknet_0_net892;
 wire clknet_1_0__leaf_net892;
 wire clknet_1_1__leaf_net892;
 wire clknet_0_net876;
 wire clknet_1_0__leaf_net876;
 wire clknet_1_1__leaf_net876;
 wire clknet_0_net534;
 wire clknet_1_0__leaf_net534;
 wire clknet_1_1__leaf_net534;
 wire clknet_0_net645;
 wire clknet_1_0__leaf_net645;
 wire clknet_1_1__leaf_net645;
 wire clknet_0_net629;
 wire clknet_1_0__leaf_net629;
 wire clknet_1_1__leaf_net629;
 wire clknet_0_net639;
 wire clknet_1_0__leaf_net639;
 wire clknet_1_1__leaf_net639;
 wire clknet_0_net641;
 wire clknet_1_0__leaf_net641;
 wire clknet_1_1__leaf_net641;
 wire clknet_0_net533;
 wire clknet_1_0__leaf_net533;
 wire clknet_1_1__leaf_net533;
 wire clknet_0_net556;
 wire clknet_1_0__leaf_net556;
 wire clknet_1_1__leaf_net556;
 wire clknet_0_net649;
 wire clknet_1_0__leaf_net649;
 wire clknet_1_1__leaf_net649;
 wire clknet_0_net540;
 wire clknet_1_0__leaf_net540;
 wire clknet_1_1__leaf_net540;
 wire clknet_0_net532;
 wire clknet_1_0__leaf_net532;
 wire clknet_1_1__leaf_net532;
 wire clknet_0_net967;
 wire clknet_1_0__leaf_net967;
 wire clknet_1_1__leaf_net967;
 wire clknet_0_net562;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_1__leaf_net562;
 wire clknet_0_net679;
 wire clknet_1_0__leaf_net679;
 wire clknet_1_1__leaf_net679;
 wire clknet_0_net674;
 wire clknet_1_0__leaf_net674;
 wire clknet_1_1__leaf_net674;
 wire clknet_0_net574;
 wire clknet_1_0__leaf_net574;
 wire clknet_1_1__leaf_net574;
 wire clknet_0_net578;
 wire clknet_1_0__leaf_net578;
 wire clknet_1_1__leaf_net578;
 wire clknet_0_net821;
 wire clknet_1_0__leaf_net821;
 wire clknet_1_1__leaf_net821;
 wire clknet_0_net440;
 wire clknet_1_0__leaf_net440;
 wire clknet_1_1__leaf_net440;
 wire clknet_0_net441;
 wire clknet_1_0__leaf_net441;
 wire clknet_1_1__leaf_net441;
 wire clknet_0_net584;
 wire clknet_1_0__leaf_net584;
 wire clknet_1_1__leaf_net584;
 wire clknet_0_net972;
 wire clknet_1_0__leaf_net972;
 wire clknet_1_1__leaf_net972;
 wire clknet_0_net840;
 wire clknet_1_0__leaf_net840;
 wire clknet_1_1__leaf_net840;
 wire clknet_0_net823;
 wire clknet_1_0__leaf_net823;
 wire clknet_1_1__leaf_net823;
 wire clknet_0_net83;
 wire clknet_1_0__leaf_net83;
 wire clknet_1_1__leaf_net83;
 wire clknet_0_net85;
 wire clknet_1_0__leaf_net85;
 wire clknet_1_1__leaf_net85;
 wire clknet_0_net103;
 wire clknet_1_0__leaf_net103;
 wire clknet_1_1__leaf_net103;
 wire clknet_0_net365;
 wire clknet_1_0__leaf_net365;
 wire clknet_1_1__leaf_net365;
 wire clknet_0_net370;
 wire clknet_1_0__leaf_net370;
 wire clknet_1_1__leaf_net370;
 wire clknet_0_net367;
 wire clknet_1_0__leaf_net367;
 wire clknet_1_1__leaf_net367;
 wire clknet_0_net81;
 wire clknet_1_0__leaf_net81;
 wire clknet_1_1__leaf_net81;
 wire clknet_0_net339;
 wire clknet_1_0__leaf_net339;
 wire clknet_1_1__leaf_net339;
 wire clknet_0_net210;
 wire clknet_1_0__leaf_net210;
 wire clknet_1_1__leaf_net210;
 wire clknet_0_net78;
 wire clknet_1_0__leaf_net78;
 wire clknet_1_1__leaf_net78;
 wire clknet_0_net346;
 wire clknet_1_0__leaf_net346;
 wire clknet_1_1__leaf_net346;
 wire clknet_0_net478;
 wire clknet_1_0__leaf_net478;
 wire clknet_1_1__leaf_net478;
 wire clknet_0_net201;
 wire clknet_1_0__leaf_net201;
 wire clknet_1_1__leaf_net201;
 wire clknet_0_net471;
 wire clknet_1_0__leaf_net471;
 wire clknet_1_1__leaf_net471;
 wire clknet_0_net89;
 wire clknet_1_0__leaf_net89;
 wire clknet_1_1__leaf_net89;
 wire clknet_0_net364;
 wire clknet_1_0__leaf_net364;
 wire clknet_1_1__leaf_net364;
 wire clknet_0_net501;
 wire clknet_1_0__leaf_net501;
 wire clknet_1_1__leaf_net501;
 wire clknet_0_net225;
 wire clknet_1_0__leaf_net225;
 wire clknet_1_1__leaf_net225;
 wire clknet_0_net227;
 wire clknet_1_0__leaf_net227;
 wire clknet_1_1__leaf_net227;
 wire net213;
 wire net231;
 wire net408;
 wire net661;
 wire net970;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;

 sky130_fd_sc_hd__nand3_2 c100 (.A(net67),
    .B(net71),
    .C(net997),
    .Y(net75));
 sky130_fd_sc_hd__and3_1 c101 (.A(net72),
    .B(net70),
    .C(net18),
    .X(net76));
 sky130_fd_sc_hd__nand3b_4 c102 (.A_N(net64),
    .B(net986),
    .C(net71),
    .Y(net77));
 sky130_fd_sc_hd__buf_4 c103 (.A(clknet_1_0__leaf_net823),
    .X(net78));
 sky130_fd_sc_hd__inv_6 c232_13 (.A(clknet_1_0__leaf_net913),
    .Y(net1021));
 sky130_fd_sc_hd__or4bb_2 c105 (.A(net70),
    .B(net28),
    .C_N(net74),
    .D_N(net68),
    .X(net79));
 sky130_fd_sc_hd__o2111ai_1 c106 (.A1(net66),
    .A2(net76),
    .B1(net69),
    .C1(net46),
    .D1(net979),
    .Y(net80));
 sky130_fd_sc_hd__or2_1 c107 (.A(net74),
    .B(clknet_1_0__leaf_net823),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net54),
    .A1(net986),
    .A2(net72),
    .A3(net29),
    .S0(net979),
    .S1(net1004),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net67),
    .A1(net72),
    .A2(net1020),
    .A3(net993),
    .S0(clknet_1_0__leaf_net78),
    .S1(clknet_1_0__leaf_net823),
    .X(net83));
 sky130_fd_sc_hd__nand2_1 c110 (.A(net18),
    .B(net947),
    .Y(net84));
 sky130_fd_sc_hd__and3b_4 c111 (.A_N(net75),
    .B(clknet_1_1__leaf_net83),
    .C(net983),
    .X(net85));
 sky130_fd_sc_hd__and3_1 c112 (.A(net947),
    .B(net84),
    .C(net968),
    .X(net86));
 sky130_fd_sc_hd__inv_1 c113 (.A(net756),
    .Y(net87));
 sky130_fd_sc_hd__nand2_2 c114 (.A(net939),
    .B(net52),
    .Y(net88));
 sky130_fd_sc_hd__nor3b_1 c115 (.A(clknet_1_0__leaf_net78),
    .B(net84),
    .C_N(net87),
    .Y(net89));
 sky130_fd_sc_hd__dfbbn_1 c116 (.CLK_N(clknet_4_10_0_clk),
    .D(net1050),
    .RESET_B(net61),
    .SET_B(net88),
    .Q(net91),
    .Q_N(net90));
 sky130_fd_sc_hd__inv_6 c117 (.A(net757),
    .Y(net92));
 sky130_fd_sc_hd__or3_1 c118 (.A(net986),
    .B(net934),
    .C(net86),
    .X(net93));
 sky130_fd_sc_hd__sdfbbn_1 c119 (.CLK_N(clknet_4_10_0_clk),
    .D(net938),
    .RESET_B(net93),
    .SCD(net88),
    .SCE(net979),
    .SET_B(net92),
    .Q(net95),
    .Q_N(net94));
 sky130_fd_sc_hd__sdfrbp_1 c120 (.CLK(clknet_4_10_0_clk),
    .D(net95),
    .RESET_B(net73),
    .SCD(net997),
    .SCE(net92),
    .Q(net97),
    .Q_N(net96));
 sky130_fd_sc_hd__sdfrbp_1 c121 (.CLK(clknet_4_10_0_clk),
    .D(net28),
    .RESET_B(net92),
    .SCD(net88),
    .SCE(net937),
    .Q(net99),
    .Q_N(net98));
 sky130_fd_sc_hd__and3b_1 c122 (.A_N(net99),
    .B(net94),
    .C(net92),
    .X(net100));
 sky130_fd_sc_hd__nand3_2 c123 (.A(net93),
    .B(net87),
    .C(net61),
    .Y(net101));
 sky130_fd_sc_hd__or4bb_1 c124 (.A(net93),
    .B(net90),
    .C_N(net974),
    .D_N(net101),
    .X(net102));
 sky130_fd_sc_hd__and3_4 c125 (.A(net72),
    .B(clknet_1_0__leaf_net85),
    .C(net92),
    .X(net103));
 sky130_fd_sc_hd__nand2b_4 c126 (.A_N(net92),
    .B(net101),
    .Y(net104));
 sky130_fd_sc_hd__or3_4 c127 (.A(net52),
    .B(net100),
    .C(net104),
    .X(net105));
 sky130_fd_sc_hd__sdfbbp_1 c128 (.CLK(clknet_4_10_0_clk),
    .D(clknet_1_0__leaf_net103),
    .RESET_B(net105),
    .SCD(net1057),
    .SCE(net104),
    .SET_B(net92),
    .Q(net107),
    .Q_N(net106));
 sky130_fd_sc_hd__mux4_4 c129 (.A0(net48),
    .A1(net88),
    .A2(net98),
    .A3(net86),
    .S0(net105),
    .S1(net791),
    .X(net108));
 sky130_fd_sc_hd__mux4_4 c130 (.A0(net107),
    .A1(clknet_1_1__leaf_net103),
    .A2(net105),
    .A3(net87),
    .S0(net104),
    .S1(net835),
    .X(net109));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net106),
    .A1(net105),
    .A2(net104),
    .A3(net87),
    .S0(net790),
    .S1(net835),
    .X(net110));
 sky130_fd_sc_hd__or2b_1 c132 (.A(net928),
    .B_N(net929),
    .X(net111));
 sky130_fd_sc_hd__nor2b_4 c133 (.A(net942),
    .B_N(net927),
    .Y(net112));
 sky130_fd_sc_hd__nand2b_4 c134 (.A_N(net943),
    .B(net937),
    .Y(net113));
 sky130_fd_sc_hd__nor2b_4 c135 (.A(net945),
    .B_N(net1006),
    .Y(net114));
 sky130_fd_sc_hd__nor2_8 c136 (.A(net947),
    .B(net1006),
    .Y(net115));
 sky130_fd_sc_hd__or2b_4 c137 (.A(net924),
    .B_N(net115),
    .X(net116));
 sky130_fd_sc_hd__and2_2 c138 (.A(net923),
    .B(net111),
    .X(net117));
 sky130_fd_sc_hd__nand2_1 c139 (.A(net117),
    .B(net116),
    .Y(net118));
 sky130_fd_sc_hd__nand2_1 c140 (.A(net118),
    .B(net929),
    .Y(net119));
 sky130_fd_sc_hd__nor2_4 c141 (.A(net117),
    .B(net114),
    .Y(net120));
 sky130_fd_sc_hd__or2b_4 c142 (.A(net116),
    .B_N(net111),
    .X(net121));
 sky130_fd_sc_hd__nor2b_2 c143 (.A(net115),
    .B_N(net120),
    .Y(net122));
 sky130_fd_sc_hd__or2_4 c144 (.A(net111),
    .B(net932),
    .X(net123));
 sky130_fd_sc_hd__or3_4 c145 (.A(net123),
    .B(net1006),
    .C(net120),
    .X(net124));
 sky130_fd_sc_hd__or2_2 c146 (.A(net932),
    .B(net119),
    .X(net125));
 sky130_fd_sc_hd__nand2_2 c147 (.A(net122),
    .B(net118),
    .Y(net126));
 sky130_fd_sc_hd__nor3_4 c148 (.A(net119),
    .B(net943),
    .C(net1006),
    .Y(net127));
 sky130_fd_sc_hd__a2111oi_4 c149 (.A1(net127),
    .A2(net120),
    .B1(net124),
    .C1(net1006),
    .D1(net121),
    .Y(net128));
 sky130_fd_sc_hd__or2_4 c150 (.A(net119),
    .B(net122),
    .X(net129));
 sky130_fd_sc_hd__mux4_1 c151 (.A0(net116),
    .A1(net126),
    .A2(net129),
    .A3(net124),
    .S0(net1038),
    .S1(net112),
    .X(net130));
 sky130_fd_sc_hd__or4bb_4 c152 (.A(net120),
    .B(net130),
    .C_N(net996),
    .D_N(net1038),
    .X(net131));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net130),
    .A1(net125),
    .A2(net123),
    .A3(net131),
    .S0(net928),
    .S1(net112),
    .X(net132));
 sky130_fd_sc_hd__nand3_2 c154 (.A(net16),
    .B(net122),
    .C(net129),
    .Y(net133));
 sky130_fd_sc_hd__nor2b_1 c155 (.A(net122),
    .B_N(net133),
    .Y(net134));
 sky130_fd_sc_hd__nor2b_1 c156 (.A(net125),
    .B_N(net134),
    .Y(net135));
 sky130_fd_sc_hd__nand2_1 c157 (.A(net4),
    .B(net14),
    .Y(net136));
 sky130_fd_sc_hd__and2_1 c158 (.A(net132),
    .B(net136),
    .X(net137));
 sky130_fd_sc_hd__nor2_2 c159 (.A(net129),
    .B(net124),
    .Y(net138));
 sky130_fd_sc_hd__nor2_8 c160 (.A(net15),
    .B(net129),
    .Y(net139));
 sky130_fd_sc_hd__nand3_2 c161 (.A(net925),
    .B(net136),
    .C(net135),
    .Y(net140));
 sky130_fd_sc_hd__and2_1 c162 (.A(net17),
    .B(net135),
    .X(net141));
 sky130_fd_sc_hd__nand2_4 c163 (.A(net140),
    .B(net139),
    .Y(net142));
 sky130_fd_sc_hd__nor2b_4 c164 (.A(net138),
    .B_N(net139),
    .Y(net143));
 sky130_fd_sc_hd__nor2_1 c165 (.A(net136),
    .B(net117),
    .Y(net144));
 sky130_fd_sc_hd__nand2b_1 c166 (.A_N(net135),
    .B(net132),
    .Y(net145));
 sky130_fd_sc_hd__mux4_2 c167 (.A0(net11),
    .A1(net926),
    .A2(net144),
    .A3(net117),
    .S0(net139),
    .S1(net944),
    .X(net146));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net10),
    .A1(net936),
    .A2(net129),
    .A3(net139),
    .S0(net998),
    .S1(net926),
    .X(net147));
 sky130_fd_sc_hd__nand3_2 c169 (.A(net998),
    .B(net138),
    .C(net143),
    .Y(net148));
 sky130_fd_sc_hd__and3_1 c170 (.A(net117),
    .B(net126),
    .C(net147),
    .X(net149));
 sky130_fd_sc_hd__nand2b_4 c171 (.A_N(net134),
    .B(net146),
    .Y(net150));
 sky130_fd_sc_hd__o2111ai_4 c172 (.A1(net144),
    .A2(net139),
    .B1(net148),
    .C1(net992),
    .D1(net985),
    .Y(net151));
 sky130_fd_sc_hd__nor3_1 c173 (.A(net138),
    .B(net117),
    .C(net985),
    .Y(net152));
 sky130_fd_sc_hd__or2_4 c174 (.A(net149),
    .B(net152),
    .X(net153));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net143),
    .A1(net927),
    .A2(net15),
    .A3(net117),
    .S0(net153),
    .S1(net947),
    .X(net154));
 sky130_fd_sc_hd__or2b_2 c176 (.A(net131),
    .B_N(net132),
    .X(net155));
 sky130_fd_sc_hd__and2_1 c177 (.A(net22),
    .B(net5),
    .X(net156));
 sky130_fd_sc_hd__and2_1 c178 (.A(net35),
    .B(net22),
    .X(net157));
 sky130_fd_sc_hd__and2b_2 c179 (.A_N(net36),
    .B(net156),
    .X(net158));
 sky130_fd_sc_hd__nor2_1 c180 (.A(net141),
    .B(net155),
    .Y(net159));
 sky130_fd_sc_hd__and2b_1 c181 (.A_N(net159),
    .B(net121),
    .X(net160));
 sky130_fd_sc_hd__nand3b_2 c182 (.A_N(net134),
    .B(net157),
    .C(net982),
    .Y(net161));
 sky130_fd_sc_hd__inv_4 c183 (.A(net809),
    .Y(net162));
 sky130_fd_sc_hd__and3_2 c184 (.A(net37),
    .B(net156),
    .C(net982),
    .X(net163));
 sky130_fd_sc_hd__or2b_1 c185 (.A(net148),
    .B_N(net162),
    .X(net164));
 sky130_fd_sc_hd__a2111oi_2 c186 (.A1(net945),
    .A2(net14),
    .B1(net155),
    .C1(net161),
    .D1(net131),
    .Y(net165));
 sky130_fd_sc_hd__sdfbbn_2 c187 (.CLK_N(clknet_4_2_0_clk),
    .D(net156),
    .RESET_B(net978),
    .SCD(net163),
    .SCE(net1004),
    .SET_B(net140),
    .Q(net167),
    .Q_N(net166));
 sky130_fd_sc_hd__or4bb_4 c188 (.A(net137),
    .B(net140),
    .C_N(net131),
    .D_N(net1007),
    .X(net168));
 sky130_fd_sc_hd__buf_1 c189 (.A(net808),
    .X(net169));
 sky130_fd_sc_hd__or4bb_1 c190 (.A(net155),
    .B(net162),
    .C_N(net168),
    .D_N(net982),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 c191 (.A0(net145),
    .A1(net37),
    .A2(net169),
    .A3(net142),
    .S0(net164),
    .S1(net163),
    .X(net171));
 sky130_fd_sc_hd__sdfbbn_1 c192 (.CLK_N(clknet_4_2_0_clk),
    .D(net169),
    .RESET_B(net156),
    .SCD(net163),
    .SCE(net945),
    .SET_B(net837),
    .Q(net173),
    .Q_N(net172));
 sky130_fd_sc_hd__and3_1 c193 (.A(net170),
    .B(net169),
    .C(net837),
    .X(net174));
 sky130_fd_sc_hd__buf_6 c194 (.A(net828),
    .X(net175));
 sky130_fd_sc_hd__mux4_4 c195 (.A0(net32),
    .A1(net170),
    .A2(net131),
    .A3(net163),
    .S0(net947),
    .S1(net837),
    .X(net176));
 sky130_fd_sc_hd__or4bb_1 c196 (.A(net163),
    .B(net145),
    .C_N(net172),
    .D_N(net1002),
    .X(net177));
 sky130_fd_sc_hd__or4bb_1 c197 (.A(net175),
    .B(net169),
    .C_N(net809),
    .D_N(net1002),
    .X(net178));
 sky130_fd_sc_hd__or3_4 c198 (.A(net40),
    .B(net29),
    .C(net1004),
    .X(net179));
 sky130_fd_sc_hd__and2_1 c199 (.A(net52),
    .B(net43),
    .X(net180));
 sky130_fd_sc_hd__and2b_1 c200 (.A_N(net154),
    .B(net36),
    .X(net181));
 sky130_fd_sc_hd__nor2_1 c201 (.A(net54),
    .B(net154),
    .Y(net182));
 sky130_fd_sc_hd__and2_0 c202 (.A(net51),
    .B(net2),
    .X(net183));
 sky130_fd_sc_hd__buf_1 c203 (.A(net738),
    .X(net184));
 sky130_fd_sc_hd__or2_1 c204 (.A(net184),
    .B(net968),
    .X(net185));
 sky130_fd_sc_hd__nor2b_1 c205 (.A(net164),
    .B_N(net43),
    .Y(net186));
 sky130_fd_sc_hd__nor2_1 c206 (.A(net175),
    .B(net43),
    .Y(net187));
 sky130_fd_sc_hd__or3b_1 c207 (.A(net186),
    .B(net54),
    .C_N(net52),
    .X(net188));
 sky130_fd_sc_hd__or4bb_1 c208 (.A(net162),
    .B(net184),
    .C_N(net187),
    .D_N(net1008),
    .X(net189));
 sky130_fd_sc_hd__inv_4 c209 (.A(net738),
    .Y(net190));
 sky130_fd_sc_hd__nor2_2 c210 (.A(net149),
    .B(net947),
    .Y(net191));
 sky130_fd_sc_hd__inv_8 c211 (.A(net803),
    .Y(net192));
 sky130_fd_sc_hd__and2_1 c212 (.A(net175),
    .B(net54),
    .X(net193));
 sky130_fd_sc_hd__nand2b_1 c213 (.A_N(net159),
    .B(net988),
    .Y(net194));
 sky130_fd_sc_hd__nor2b_2 c214 (.A(net182),
    .B_N(net193),
    .Y(net195));
 sky130_fd_sc_hd__and2b_1 c215 (.A_N(net189),
    .B(net187),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 c216 (.A(net803),
    .X(net197));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net194),
    .A1(net157),
    .A2(net193),
    .A3(net924),
    .S0(net166),
    .S1(net185),
    .X(net198));
 sky130_fd_sc_hd__nand2_1 c218 (.A(net185),
    .B(net168),
    .Y(net199));
 sky130_fd_sc_hd__and2b_4 c219 (.A_N(net199),
    .B(net185),
    .X(net200));
 sky130_fd_sc_hd__or3_4 c220 (.A(clknet_1_1__leaf_net78),
    .B(net985),
    .C(net160),
    .X(net201));
 sky130_fd_sc_hd__buf_1 c221 (.A(net915),
    .X(net202));
 sky130_fd_sc_hd__nand2b_1 c222 (.A_N(net202),
    .B(net187),
    .Y(net203));
 sky130_fd_sc_hd__inv_12 c223 (.A(net741),
    .Y(net204));
 sky130_fd_sc_hd__clkbuf_1 c224 (.A(net803),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 c225 (.A(net741),
    .X(net206));
 sky130_fd_sc_hd__or4bb_2 c226 (.A(net206),
    .B(clknet_1_1__leaf_net78),
    .C_N(net139),
    .D_N(net202),
    .X(net207));
 sky130_fd_sc_hd__a2111o_2 c227 (.A1(net1004),
    .A2(net143),
    .B1(net197),
    .C1(net139),
    .D1(net204),
    .X(net208));
 sky130_fd_sc_hd__and3_1 c228 (.A(net160),
    .B(net202),
    .C(net833),
    .X(net209));
 sky130_fd_sc_hd__and3b_2 c229 (.A_N(net160),
    .B(clknet_1_1__leaf_net81),
    .C(net75),
    .X(net210));
 sky130_fd_sc_hd__or4bb_1 c230 (.A(net205),
    .B(net209),
    .C_N(net65),
    .D_N(net999),
    .X(net211));
 sky130_fd_sc_hd__nor3_1 c231 (.A(net43),
    .B(net927),
    .C(net197),
    .Y(net212));
 sky130_fd_sc_hd__inv_6 c250_20 (.A(clknet_1_1__leaf_net913),
    .Y(net1028));
 sky130_fd_sc_hd__nand3b_2 c233 (.A_N(net196),
    .B(net39),
    .C(net1027),
    .Y(net214));
 sky130_fd_sc_hd__nor3b_1 c234 (.A(net212),
    .B(net204),
    .C_N(net833),
    .Y(net215));
 sky130_fd_sc_hd__o2111ai_4 c235 (.A1(net203),
    .A2(net1026),
    .B1(clknet_1_1__leaf_net214),
    .C1(net987),
    .D1(net795),
    .Y(net216));
 sky130_fd_sc_hd__or4bb_1 c236 (.A(net75),
    .B(net970),
    .C_N(net979),
    .D_N(net1025),
    .X(net217));
 sky130_fd_sc_hd__mux4_4 c237 (.A0(net1024),
    .A1(clknet_1_0__leaf_net201),
    .A2(net197),
    .A3(clknet_1_0__leaf_net210),
    .S0(net204),
    .S1(clknet_1_0__leaf_net214),
    .X(net218));
 sky130_fd_sc_hd__mux4_4 c238 (.A0(net29),
    .A1(clknet_1_0__leaf_net214),
    .A2(net1023),
    .A3(net987),
    .S0(clknet_1_0__leaf_net210),
    .S1(net979),
    .X(net219));
 sky130_fd_sc_hd__mux4_2 c239 (.A0(net218),
    .A1(net77),
    .A2(clknet_1_0__leaf_net214),
    .A3(net1022),
    .S0(net970),
    .S1(clknet_1_0__leaf_net839),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net196),
    .A1(clknet_1_0__leaf_net201),
    .A2(net987),
    .A3(clknet_1_0__leaf_net210),
    .S0(net828),
    .S1(clknet_1_0__leaf_net839),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net215),
    .A1(net1021),
    .A2(clknet_1_0__leaf_net210),
    .A3(net987),
    .S0(net832),
    .S1(clknet_1_1__leaf_net839),
    .X(net222));
 sky130_fd_sc_hd__and2b_2 c242 (.A_N(net215),
    .B(clknet_1_0__leaf_net214),
    .X(net223));
 sky130_fd_sc_hd__inv_2 c243 (.A(net755),
    .Y(net224));
 sky130_fd_sc_hd__nand3_1 c244 (.A(net224),
    .B(clknet_1_0__leaf_net89),
    .C(net1008),
    .Y(net225));
 sky130_fd_sc_hd__inv_1 c245 (.A(net754),
    .Y(net226));
 sky130_fd_sc_hd__and3_1 c246 (.A(net91),
    .B(net52),
    .C(clknet_1_0__leaf_net225),
    .X(net227));
 sky130_fd_sc_hd__or2_2 c247 (.A(net97),
    .B(clknet_1_1__leaf_net223),
    .X(net228));
 sky130_fd_sc_hd__inv_1 c248 (.A(net768),
    .Y(net229));
 sky130_fd_sc_hd__nor2_2 c249 (.A(net197),
    .B(net193),
    .Y(net230));
 sky130_fd_sc_hd__nand2b_1 c25 (.A_N(net8),
    .B(net939),
    .Y(net0));
 sky130_fd_sc_hd__inv_2 c423_24 (.A(clknet_1_0__leaf_net914),
    .Y(net1032));
 sky130_fd_sc_hd__inv_2 c251 (.A(net768),
    .Y(net232));
 sky130_fd_sc_hd__inv_1 c252 (.A(net794),
    .Y(net233));
 sky130_fd_sc_hd__and2_1 c253 (.A(net1008),
    .B(net1031),
    .X(net234));
 sky130_fd_sc_hd__or4bb_4 c254 (.A(net88),
    .B(net97),
    .C_N(net230),
    .D_N(clknet_1_0__leaf_net214),
    .X(net235));
 sky130_fd_sc_hd__mux4_2 c255 (.A0(net101),
    .A1(net215),
    .A2(clknet_1_0__leaf_net227),
    .A3(net979),
    .S0(net985),
    .S1(net988),
    .X(net236));
 sky130_fd_sc_hd__a2111o_4 c256 (.A1(net86),
    .A2(net924),
    .B1(net48),
    .C1(net797),
    .D1(clknet_1_1__leaf_net840),
    .X(net237));
 sky130_fd_sc_hd__or3b_2 c257 (.A(net61),
    .B(net1008),
    .C_N(net988),
    .X(net238));
 sky130_fd_sc_hd__and3b_2 c258 (.A_N(net226),
    .B(net233),
    .C(clknet_1_0__leaf_net840),
    .X(net239));
 sky130_fd_sc_hd__or3b_4 c259 (.A(net1030),
    .B(net238),
    .C_N(clknet_1_0__leaf_net840),
    .X(net240));
 sky130_fd_sc_hd__and2_2 c26 (.A(net0),
    .B(net938),
    .X(net1));
 sky130_fd_sc_hd__or3_2 c260 (.A(net239),
    .B(clknet_1_0__leaf_net223),
    .C(net834),
    .X(net241));
 sky130_fd_sc_hd__mux4_4 c261 (.A0(net237),
    .A1(clknet_1_0__leaf_net241),
    .A2(net104),
    .A3(net979),
    .S0(net5),
    .S1(clknet_1_1__leaf_net840),
    .X(net242));
 sky130_fd_sc_hd__mux4_4 c262 (.A0(net229),
    .A1(net1029),
    .A2(clknet_1_0__leaf_net240),
    .A3(clknet_1_1__leaf_net241),
    .S0(net797),
    .S1(clknet_1_0__leaf_net840),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(clknet_1_1__leaf_net225),
    .A1(clknet_1_0__leaf_net241),
    .A2(net75),
    .A3(net947),
    .S0(net79),
    .S1(net797),
    .X(net244));
 sky130_fd_sc_hd__nand3_1 c264 (.A(net115),
    .B(net946),
    .C(net1038),
    .Y(net245));
 sky130_fd_sc_hd__or2b_1 c265 (.A(net125),
    .B_N(net131),
    .X(net246));
 sky130_fd_sc_hd__or2b_1 c266 (.A(net1038),
    .B_N(net928),
    .X(net247));
 sky130_fd_sc_hd__and2b_2 c267 (.A_N(net944),
    .B(net995),
    .X(net248));
 sky130_fd_sc_hd__nor2_1 c268 (.A(net946),
    .B(net248),
    .Y(net249));
 sky130_fd_sc_hd__nand3b_1 c269 (.A_N(net247),
    .B(net115),
    .C(net1063),
    .Y(net250));
 sky130_fd_sc_hd__and2_4 c27 (.A(net944),
    .B(net936),
    .X(net2));
 sky130_fd_sc_hd__or4bb_4 c270 (.A(net995),
    .B(net114),
    .C_N(net248),
    .D_N(net1038),
    .X(net251));
 sky130_fd_sc_hd__nand2_4 c271 (.A(net251),
    .B(net929),
    .Y(net252));
 sky130_fd_sc_hd__or2_2 c272 (.A(net249),
    .B(net123),
    .X(net253));
 sky130_fd_sc_hd__and2_4 c273 (.A(net248),
    .B(net245),
    .X(net254));
 sky130_fd_sc_hd__and2_1 c274 (.A(net114),
    .B(net247),
    .X(net255));
 sky130_fd_sc_hd__and2_1 c275 (.A(net252),
    .B(net131),
    .X(net256));
 sky130_fd_sc_hd__a2111o_1 c276 (.A1(net253),
    .A2(net256),
    .B1(net254),
    .C1(net115),
    .D1(net1063),
    .X(net257));
 sky130_fd_sc_hd__and2_1 c277 (.A(net929),
    .B(net248),
    .X(net258));
 sky130_fd_sc_hd__nor3b_1 c278 (.A(net256),
    .B(net1062),
    .C_N(net252),
    .Y(net259));
 sky130_fd_sc_hd__or2_4 c279 (.A(net248),
    .B(net255),
    .X(net260));
 sky130_fd_sc_hd__or2b_2 c28 (.A(net931),
    .B_N(net940),
    .X(net3));
 sky130_fd_sc_hd__nor2b_2 c280 (.A(net257),
    .B_N(net132),
    .Y(net261));
 sky130_fd_sc_hd__nand2b_1 c281 (.A_N(net131),
    .B(net251),
    .Y(net262));
 sky130_fd_sc_hd__nand3_1 c282 (.A(net262),
    .B(net257),
    .C(net261),
    .Y(net959));
 sky130_fd_sc_hd__and2_1 c283 (.A(net245),
    .B(net258),
    .X(net263));
 sky130_fd_sc_hd__mux4_2 c284 (.A0(net250),
    .A1(net263),
    .A2(net249),
    .A3(net1063),
    .S0(net254),
    .S1(net261),
    .X(net264));
 sky130_fd_sc_hd__o2111ai_1 c285 (.A1(net258),
    .A2(net114),
    .B1(net264),
    .C1(net261),
    .D1(net981),
    .Y(net265));
 sky130_fd_sc_hd__nand2_1 c286 (.A(net148),
    .B(net152),
    .Y(net266));
 sky130_fd_sc_hd__nor3b_1 c287 (.A(net8),
    .B(net266),
    .C_N(net143),
    .Y(net267));
 sky130_fd_sc_hd__and3b_1 c288 (.A_N(net135),
    .B(net985),
    .C(net924),
    .X(net268));
 sky130_fd_sc_hd__and3b_2 c289 (.A_N(net266),
    .B(net135),
    .C(net985),
    .X(net269));
 sky130_fd_sc_hd__nor2_1 c29 (.A(net926),
    .B(net1),
    .Y(net4));
 sky130_fd_sc_hd__and3_1 c290 (.A(net261),
    .B(net153),
    .C(net269),
    .X(net270));
 sky130_fd_sc_hd__and3_1 c291 (.A(net267),
    .B(net125),
    .C(net253),
    .X(net271));
 sky130_fd_sc_hd__nor2_1 c292 (.A(net254),
    .B(net262),
    .Y(net272));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(net13),
    .A1(net271),
    .A2(net270),
    .A3(net17),
    .S0(net8),
    .S1(net985),
    .X(net273));
 sky130_fd_sc_hd__and2_2 c294 (.A(net259),
    .B(net153),
    .X(net274));
 sky130_fd_sc_hd__mux4_4 c295 (.A0(net273),
    .A1(net925),
    .A2(net259),
    .A3(net270),
    .S0(net936),
    .S1(net981),
    .X(net275));
 sky130_fd_sc_hd__mux4_4 c296 (.A0(net262),
    .A1(net273),
    .A2(net259),
    .A3(net154),
    .S0(net985),
    .S1(net125),
    .X(net276));
 sky130_fd_sc_hd__and3_1 c297 (.A(net151),
    .B(net269),
    .C(net268),
    .X(net277));
 sky130_fd_sc_hd__and3b_1 c298 (.A_N(net270),
    .B(net269),
    .C(net810),
    .X(net278));
 sky130_fd_sc_hd__and2_2 c299 (.A(net261),
    .B(net810),
    .X(net279));
 sky130_fd_sc_hd__nor2b_2 c30 (.A(net3),
    .B_N(net0),
    .Y(net5));
 sky130_fd_sc_hd__nand2_2 c300 (.A(net277),
    .B(net253),
    .Y(net280));
 sky130_fd_sc_hd__buf_1 c301 (.A(net911),
    .X(net281));
 sky130_fd_sc_hd__and3_1 c302 (.A(net936),
    .B(net267),
    .C(net810),
    .X(net282));
 sky130_fd_sc_hd__or3b_1 c303 (.A(net152),
    .B(net944),
    .C_N(net142),
    .X(net283));
 sky130_fd_sc_hd__and2b_1 c304 (.A_N(net283),
    .B(net811),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net283),
    .A1(net8),
    .A2(net280),
    .A3(net252),
    .S0(net133),
    .S1(net284),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net284),
    .A1(net259),
    .A2(net280),
    .A3(net142),
    .S0(net270),
    .S1(net844),
    .X(net286));
 sky130_fd_sc_hd__mux4_2 c307 (.A0(net268),
    .A1(net267),
    .A2(net126),
    .A3(net284),
    .S0(net845),
    .S1(net846),
    .X(net287));
 sky130_fd_sc_hd__or4bb_4 c308 (.A(net146),
    .B(net139),
    .C_N(net279),
    .D_N(net941),
    .X(net288));
 sky130_fd_sc_hd__inv_1 c309 (.Y(net289));
 sky130_fd_sc_hd__and3_1 c31 (.A(net2),
    .B(net0),
    .C(net928),
    .X(net6));
 sky130_fd_sc_hd__nor3b_2 c310 (.A(net140),
    .B(net17),
    .C_N(net1002),
    .Y(net290));
 sky130_fd_sc_hd__sdfbbp_1 c311 (.CLK(clknet_4_2_0_clk),
    .D(net161),
    .RESET_B(net288),
    .SCD(net165),
    .SCE(net2),
    .SET_B(net141),
    .Q(net292),
    .Q_N(net291));
 sky130_fd_sc_hd__buf_16 c312 (.A(net753),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 c313 (.A(net803),
    .X(net953));
 sky130_fd_sc_hd__inv_2 c314 (.A(net911),
    .Y(net294));
 sky130_fd_sc_hd__nand2b_1 c315 (.A_N(net178),
    .B(net1000),
    .Y(net295));
 sky130_fd_sc_hd__nor2b_1 c316 (.A(net293),
    .B_N(net279),
    .Y(net296));
 sky130_fd_sc_hd__buf_1 c317 (.A(net765),
    .X(net297));
 sky130_fd_sc_hd__and2_1 c318 (.A(net295),
    .B(net982),
    .X(net298));
 sky130_fd_sc_hd__sdfbbn_2 c319 (.CLK_N(clknet_4_2_0_clk),
    .D(net165),
    .RESET_B(net293),
    .SCD(net269),
    .SCE(net290),
    .SET_B(net1002),
    .Q(net300),
    .Q_N(net299));
 sky130_fd_sc_hd__and2_1 c32 (.A(net946),
    .B(net2),
    .X(net7));
 sky130_fd_sc_hd__and2_1 c320 (.A(net292),
    .B(net271),
    .X(net301));
 sky130_fd_sc_hd__inv_1 c321 (.A(net816),
    .Y(net302));
 sky130_fd_sc_hd__a2111o_1 c322 (.A1(net24),
    .A2(net163),
    .B1(net293),
    .C1(net291),
    .D1(net1002),
    .X(net303));
 sky130_fd_sc_hd__a2111o_1 c323 (.A1(net297),
    .A2(net295),
    .B1(net298),
    .C1(net299),
    .D1(net293),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(net271),
    .A1(net301),
    .A2(net293),
    .A3(net288),
    .S0(net291),
    .S1(net178),
    .X(net305));
 sky130_fd_sc_hd__sdfbbn_2 c325 (.CLK_N(clknet_4_3_0_clk),
    .D(net298),
    .RESET_B(net304),
    .SCD(net297),
    .SCE(net292),
    .SET_B(net288),
    .Q(net307),
    .Q_N(net306));
 sky130_fd_sc_hd__sdfbbp_1 c326 (.CLK(clknet_4_3_0_clk),
    .D(net288),
    .RESET_B(net298),
    .SCD(net306),
    .SCE(net811),
    .SET_B(net1040),
    .Q(net309),
    .Q_N(net308));
 sky130_fd_sc_hd__a2111o_1 c327 (.A1(net271),
    .A2(net307),
    .B1(net163),
    .C1(net292),
    .D1(net1045),
    .X(net310));
 sky130_fd_sc_hd__sdfbbn_1 c328 (.CLK_N(clknet_4_3_0_clk),
    .D(net304),
    .RESET_B(net158),
    .SCD(net298),
    .SCE(net161),
    .SET_B(net1053),
    .Q(net312),
    .Q_N(net311));
 sky130_fd_sc_hd__o2111ai_1 c329 (.A1(net311),
    .A2(net307),
    .B1(net146),
    .C1(net924),
    .D1(net814),
    .Y(net313));
 sky130_fd_sc_hd__and2b_1 c33 (.A_N(net935),
    .B(net928),
    .X(net8));
 sky130_fd_sc_hd__and2_0 c330 (.A(net302),
    .B(net274),
    .X(net314));
 sky130_fd_sc_hd__and2b_1 c331 (.A_N(net196),
    .B(net300),
    .X(net315));
 sky130_fd_sc_hd__o2111ai_2 c332 (.A1(net294),
    .A2(net300),
    .B1(net291),
    .C1(net191),
    .D1(net845),
    .Y(net316));
 sky130_fd_sc_hd__a2111oi_2 c333 (.A1(net198),
    .A2(net927),
    .B1(net46),
    .C1(net315),
    .D1(net196),
    .Y(net317));
 sky130_fd_sc_hd__nor2b_1 c334 (.A(net934),
    .B_N(net190),
    .Y(net318));
 sky130_fd_sc_hd__inv_2 c335 (.A(net759),
    .Y(net319));
 sky130_fd_sc_hd__and2_1 c336 (.A(net191),
    .B(net315),
    .X(net320));
 sky130_fd_sc_hd__nor2b_1 c337 (.A(net1044),
    .B_N(net292),
    .Y(net321));
 sky130_fd_sc_hd__nand2_4 c338 (.A(net279),
    .B(net48),
    .Y(net322));
 sky130_fd_sc_hd__nand2b_2 c339 (.A_N(net321),
    .B(net168),
    .Y(net323));
 sky130_fd_sc_hd__or2b_2 c34 (.A(net939),
    .B_N(net7),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 c340 (.A(net910),
    .X(net324));
 sky130_fd_sc_hd__or4bb_4 c341 (.A(net324),
    .B(net319),
    .C_N(net982),
    .D_N(net166),
    .X(net325));
 sky130_fd_sc_hd__a2111o_1 c342 (.A1(net183),
    .A2(net191),
    .B1(net323),
    .C1(net48),
    .D1(net325),
    .X(net326));
 sky130_fd_sc_hd__a2111o_1 c343 (.A1(net318),
    .A2(net321),
    .B1(net968),
    .C1(net279),
    .D1(net793),
    .X(net327));
 sky130_fd_sc_hd__sdfbbn_2 c344 (.CLK_N(clknet_4_9_0_clk),
    .D(net327),
    .RESET_B(net325),
    .SCD(net291),
    .SCE(net814),
    .SET_B(net1001),
    .Q(net966),
    .Q_N(net328));
 sky130_fd_sc_hd__clkbuf_1 c345 (.A(net758),
    .X(net329));
 sky130_fd_sc_hd__inv_1 c346 (.A(net765),
    .Y(net330));
 sky130_fd_sc_hd__nor2b_1 c347 (.A(net168),
    .B_N(net320),
    .Y(net331));
 sky130_fd_sc_hd__or2b_2 c348 (.A(net292),
    .B_N(net330),
    .X(net332));
 sky130_fd_sc_hd__a2111oi_1 c349 (.A1(net317),
    .A2(net55),
    .B1(net158),
    .C1(net320),
    .D1(net982),
    .Y(net333));
 sky130_fd_sc_hd__nand2_2 c35 (.A(net7),
    .B(net1),
    .Y(net10));
 sky130_fd_sc_hd__mux4_4 c350 (.A0(net331),
    .A1(net977),
    .A2(net274),
    .A3(net328),
    .S0(net190),
    .S1(net792),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net313),
    .A1(net321),
    .A2(net966),
    .A3(net331),
    .S0(net322),
    .S1(net848),
    .X(net335));
 sky130_fd_sc_hd__nor3b_1 c352 (.A(net200),
    .B(net77),
    .C_N(net209),
    .Y(net336));
 sky130_fd_sc_hd__or4bb_1 c353 (.A(net314),
    .B(net982),
    .C_N(net1000),
    .D_N(net1001),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 c354 (.A(net737),
    .X(net338));
 sky130_fd_sc_hd__nand3_1 c355 (.A(net980),
    .B(clknet_1_0__leaf_net81),
    .C(net811),
    .Y(net339));
 sky130_fd_sc_hd__nor3b_1 c356 (.A(net320),
    .B(net167),
    .C_N(net1001),
    .Y(net340));
 sky130_fd_sc_hd__and3_1 c357 (.A(net927),
    .B(net332),
    .C(net9),
    .X(net341));
 sky130_fd_sc_hd__buf_1 c358 (.A(net736),
    .X(net954));
 sky130_fd_sc_hd__or4bb_1 c359 (.A(net341),
    .B(net77),
    .C_N(net287),
    .D_N(net204),
    .X(net342));
 sky130_fd_sc_hd__nor2b_2 c36 (.A(net997),
    .B_N(net998),
    .Y(net11));
 sky130_fd_sc_hd__or3b_1 c360 (.A(net209),
    .B(net196),
    .C_N(net987),
    .X(net343));
 sky130_fd_sc_hd__inv_2 c361 (.A(net910),
    .Y(net344));
 sky130_fd_sc_hd__sdfrtn_1 c362 (.CLK_N(clknet_4_8_0_clk),
    .D(net221),
    .RESET_B(net192),
    .SCD(net343),
    .SCE(clknet_1_0__leaf_net210),
    .Q(net345));
 sky130_fd_sc_hd__nor2_2 c363 (.A(net207),
    .B(net167),
    .Y(net346));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net343),
    .A1(net340),
    .A2(net329),
    .A3(net408),
    .S0(net322),
    .S1(net1002),
    .X(net347));
 sky130_fd_sc_hd__and2b_1 c365 (.A_N(net345),
    .B(net795),
    .X(net348));
 sky130_fd_sc_hd__nand3_1 c366 (.A(net77),
    .B(net819),
    .C(net1002),
    .Y(net349));
 sky130_fd_sc_hd__sdfrtp_1 c367 (.CLK(clknet_4_9_0_clk),
    .D(net158),
    .RESET_B(net315),
    .SCD(net337),
    .SCE(net341),
    .Q(net350));
 sky130_fd_sc_hd__nor2b_1 c368 (.A(net338),
    .B_N(net818),
    .Y(net351));
 sky130_fd_sc_hd__or4bb_2 c369 (.A(net216),
    .B(net344),
    .C_N(net954),
    .D_N(clknet_1_0__leaf_net346),
    .X(net352));
 sky130_fd_sc_hd__or4bb_1 c37 (.A(net1),
    .B(net11),
    .C_N(net939),
    .D_N(net997),
    .X(net12));
 sky130_fd_sc_hd__mux4_4 c370 (.A0(net329),
    .A1(clknet_1_1__leaf_net339),
    .A2(net349),
    .A3(net314),
    .S0(clknet_1_0__leaf_net210),
    .S1(clknet_1_1__leaf_net201),
    .X(net353));
 sky130_fd_sc_hd__sdfrtp_1 c371 (.CLK(clknet_4_9_0_clk),
    .D(net348),
    .RESET_B(clknet_1_1__leaf_net81),
    .SCD(net287),
    .SCE(net1056),
    .Q(net354));
 sky130_fd_sc_hd__and3_2 c372 (.A(net187),
    .B(net349),
    .C(net354),
    .X(net355));
 sky130_fd_sc_hd__mux4_2 c373 (.A0(net354),
    .A1(net55),
    .A2(net355),
    .A3(net192),
    .S0(net1002),
    .S1(net850),
    .X(net356));
 sky130_fd_sc_hd__a2111o_1 c374 (.A1(net315),
    .A2(net233),
    .B1(clknet_1_0__leaf_net222),
    .C1(net230),
    .D1(net200),
    .X(net357));
 sky130_fd_sc_hd__sdfbbp_1 c375 (.CLK(clknet_4_11_0_clk),
    .D(clknet_1_1__leaf_net227),
    .RESET_B(net966),
    .SCD(clknet_1_1__leaf_net214),
    .SCE(net983),
    .SET_B(clknet_1_0__leaf_net840),
    .Q(net359),
    .Q_N(net358));
 sky130_fd_sc_hd__sdfrtp_1 c376 (.CLK(clknet_4_11_0_clk),
    .D(clknet_1_0__leaf_net240),
    .RESET_B(net988),
    .SCD(clknet_1_0__leaf_net222),
    .SCE(net1019),
    .Q(net360));
 sky130_fd_sc_hd__or4bb_1 c377 (.A(net48),
    .B(net238),
    .C_N(net104),
    .D_N(net1001),
    .X(net361));
 sky130_fd_sc_hd__a2111o_4 c378 (.A1(clknet_1_0__leaf_net352),
    .A2(net359),
    .B1(net355),
    .C1(net983),
    .D1(net1001),
    .X(net362));
 sky130_fd_sc_hd__mux4_4 c379 (.A0(net238),
    .A1(clknet_1_1__leaf_net89),
    .A2(net1018),
    .A3(net350),
    .S0(net361),
    .S1(net792),
    .X(net363));
 sky130_fd_sc_hd__nand3b_4 c38 (.A_N(net12),
    .B(net3),
    .C(net10),
    .Y(net968));
 sky130_fd_sc_hd__or4bb_1 c380 (.A(clknet_1_0__leaf_net89),
    .B(net351),
    .C_N(net360),
    .D_N(net1000),
    .X(net364));
 sky130_fd_sc_hd__or4bb_2 c381 (.A(net153),
    .B(net358),
    .C_N(net360),
    .D_N(net1017),
    .X(net365));
 sky130_fd_sc_hd__or4bb_2 c382 (.A(net232),
    .B(clknet_1_0__leaf_net365),
    .C_N(net980),
    .D_N(net983),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c383 (.A0(net238),
    .A1(clknet_1_0__leaf_net365),
    .A2(net983),
    .A3(net835),
    .S0(net836),
    .S1(net844),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c384 (.A0(clknet_1_1__leaf_net240),
    .A1(net999),
    .A2(net358),
    .A3(clknet_1_1__leaf_net365),
    .S0(net287),
    .S1(net836),
    .X(net368));
 sky130_fd_sc_hd__mux4_4 c385 (.A0(clknet_1_1__leaf_net85),
    .A1(net366),
    .A2(clknet_1_0__leaf_net364),
    .A3(net355),
    .S0(clknet_1_0__leaf_net365),
    .S1(net924),
    .X(net369));
 sky130_fd_sc_hd__mux4_4 c386 (.A0(net1016),
    .A1(clknet_1_0__leaf_net365),
    .A2(clknet_1_1__leaf_net201),
    .A3(net799),
    .S0(net844),
    .S1(net852),
    .X(net370));
 sky130_fd_sc_hd__mux4_4 c387 (.A0(clknet_1_1__leaf_net370),
    .A1(net104),
    .A2(clknet_1_1__leaf_net234),
    .A3(net798),
    .S0(net836),
    .S1(net853),
    .X(net371));
 sky130_fd_sc_hd__mux4_4 c388 (.A0(net359),
    .A1(net238),
    .A2(clknet_1_0__leaf_net364),
    .A3(clknet_1_1__leaf_net367),
    .S0(clknet_1_1__leaf_net840),
    .S1(net852),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 c389 (.A0(clknet_1_0__leaf_net367),
    .A1(net345),
    .A2(clknet_1_0__leaf_net365),
    .A3(clknet_1_0__leaf_net364),
    .S0(net842),
    .S1(net853),
    .X(net373));
 sky130_fd_sc_hd__and2_1 c39 (.A(net1054),
    .B(net11),
    .X(net13));
 sky130_fd_sc_hd__mux4_4 c390 (.A0(net373),
    .A1(net372),
    .A2(clknet_1_1__leaf_net352),
    .A3(net1015),
    .S0(clknet_1_1__leaf_net370),
    .S1(clknet_1_1__leaf_net840),
    .X(net374));
 sky130_fd_sc_hd__mux4_4 c391 (.A0(clknet_1_0__leaf_net234),
    .A1(clknet_1_1__leaf_net222),
    .A2(net924),
    .A3(net238),
    .S0(net836),
    .S1(net855),
    .X(net375));
 sky130_fd_sc_hd__sdfbbn_1 c392 (.CLK_N(clknet_4_14_0_clk),
    .D(net322),
    .RESET_B(net834),
    .SCD(net851),
    .SCE(net855),
    .SET_B(net856),
    .Q(net377),
    .Q_N(net376));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net360),
    .A1(clknet_1_0__leaf_net370),
    .A2(net989),
    .A3(clknet_1_1__leaf_net365),
    .S0(net105),
    .S1(net854),
    .X(net378));
 sky130_fd_sc_hd__sdfbbn_1 c394 (.CLK_N(clknet_4_14_0_clk),
    .D(net363),
    .RESET_B(clknet_1_1__leaf_net370),
    .SCD(net853),
    .SCE(net855),
    .SET_B(net857),
    .Q(net379));
 sky130_fd_sc_hd__mux4_2 c395 (.A0(clknet_1_1__leaf_net214),
    .A1(net361),
    .A2(net379),
    .A3(clknet_1_0__leaf_net370),
    .S0(net153),
    .S1(net376),
    .X(net380));
 sky130_fd_sc_hd__nor2b_2 c396 (.A(net261),
    .B_N(net941),
    .Y(net381));
 sky130_fd_sc_hd__or2b_1 c397 (.A(net250),
    .B_N(net381),
    .X(net382));
 sky130_fd_sc_hd__nand2_1 c398 (.A(net981),
    .B(net263),
    .Y(net383));
 sky130_fd_sc_hd__buf_16 c399 (.A(net824),
    .X(net384));
 sky130_fd_sc_hd__or4bb_2 c40 (.A(net3),
    .B(net4),
    .C_N(net8),
    .D_N(net997),
    .X(net14));
 sky130_fd_sc_hd__or2_1 c400 (.A(net263),
    .B(net261),
    .X(net385));
 sky130_fd_sc_hd__or2_2 c401 (.A(net121),
    .B(net264),
    .X(net386));
 sky130_fd_sc_hd__inv_2 c402 (.A(net824),
    .Y(net387));
 sky130_fd_sc_hd__buf_1 c403 (.A(net760),
    .X(net388));
 sky130_fd_sc_hd__clkinv_2 c404 (.A(net829),
    .Y(net389));
 sky130_fd_sc_hd__nor2b_1 c405 (.A(net384),
    .B_N(net250),
    .Y(net390));
 sky130_fd_sc_hd__nand2b_1 c406 (.A_N(net123),
    .B(net996),
    .Y(net391));
 sky130_fd_sc_hd__or2_2 c407 (.A(net387),
    .B(net389),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 c408 (.A(net760),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 c409 (.A(net769),
    .X(net394));
 sky130_fd_sc_hd__nand2b_4 c41 (.A_N(net13),
    .B(net11),
    .Y(net15));
 sky130_fd_sc_hd__nand2b_1 c410 (.A_N(net394),
    .B(net263),
    .Y(net395));
 sky130_fd_sc_hd__inv_1 c411 (.A(net776),
    .Y(net396));
 sky130_fd_sc_hd__or2b_2 c412 (.A(net392),
    .B_N(net396),
    .X(net397));
 sky130_fd_sc_hd__and3b_1 c413 (.A_N(net395),
    .B(net126),
    .C(net393),
    .X(net398));
 sky130_fd_sc_hd__inv_4 c414 (.A(net776),
    .Y(net399));
 sky130_fd_sc_hd__nor3_1 c415 (.A(net396),
    .B(net391),
    .C(net252),
    .Y(net400));
 sky130_fd_sc_hd__o2111ai_4 c416 (.A1(net400),
    .A2(net390),
    .B1(net397),
    .C1(net398),
    .D1(net387),
    .Y(net401));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net390),
    .A1(net394),
    .A2(net395),
    .A3(net401),
    .S0(net397),
    .S1(net383),
    .X(net402));
 sky130_fd_sc_hd__nand2_4 c418 (.A(net252),
    .B(net274),
    .Y(net403));
 sky130_fd_sc_hd__nand2_4 c419 (.A(net397),
    .B(net154),
    .Y(net404));
 sky130_fd_sc_hd__a2111oi_4 c42 (.A1(net7),
    .A2(net13),
    .B1(net15),
    .C1(net997),
    .D1(net2),
    .Y(net16));
 sky130_fd_sc_hd__inv_1 c420 (.A(net813),
    .Y(net405));
 sky130_fd_sc_hd__nand3_1 c421 (.A(net381),
    .B(net252),
    .C(net403),
    .Y(net406));
 sky130_fd_sc_hd__and3b_2 c422 (.A_N(net141),
    .B(net399),
    .C(net404),
    .X(net407));
 sky130_fd_sc_hd__clkinv_4 c694_25 (.A(clknet_1_1__leaf_net914),
    .Y(net1033));
 sky130_fd_sc_hd__buf_6 c424 (.A(clknet_1_0__leaf_net912),
    .X(net409));
 sky130_fd_sc_hd__or3_1 c425 (.A(net126),
    .B(net269),
    .C(net282),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 c426 (.A(net787),
    .X(net411));
 sky130_fd_sc_hd__buf_1 c427 (.A(net921),
    .X(net412));
 sky130_fd_sc_hd__or3b_1 c428 (.A(net412),
    .B(net397),
    .C_N(net281),
    .X(net413));
 sky130_fd_sc_hd__inv_1 c429 (.A(net813),
    .Y(net414));
 sky130_fd_sc_hd__mux4_2 c43 (.A0(net10),
    .A1(net931),
    .A2(net937),
    .A3(net15),
    .S0(net1),
    .S1(net16),
    .X(net17));
 sky130_fd_sc_hd__nor3_1 c430 (.A(net411),
    .B(net414),
    .C(net412),
    .Y(net415));
 sky130_fd_sc_hd__buf_1 c431 (.A(net921),
    .X(net416));
 sky130_fd_sc_hd__inv_6 c432 (.A(net922),
    .Y(net417));
 sky130_fd_sc_hd__nand3b_1 c433 (.A_N(net416),
    .B(net417),
    .C(net274),
    .Y(net418));
 sky130_fd_sc_hd__nand3_2 c434 (.A(net414),
    .B(net389),
    .C(net416),
    .Y(net419));
 sky130_fd_sc_hd__or3b_1 c435 (.A(net416),
    .B(net419),
    .C_N(clknet_1_0__leaf_net409),
    .X(net420));
 sky130_fd_sc_hd__inv_4 c436 (.A(net786),
    .Y(net421));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net417),
    .A1(net261),
    .A2(net413),
    .A3(net416),
    .S0(net661),
    .S1(net403),
    .X(net422));
 sky130_fd_sc_hd__and3_2 c438 (.A(net418),
    .B(net421),
    .C(net416),
    .X(net423));
 sky130_fd_sc_hd__mux4_4 c439 (.A0(net281),
    .A1(net417),
    .A2(net401),
    .A3(clknet_1_0__leaf_net420),
    .S0(net280),
    .S1(net975),
    .X(net424));
 sky130_fd_sc_hd__and2_1 c44 (.A(net930),
    .B(net928),
    .X(net18));
 sky130_fd_sc_hd__nand2b_1 c440 (.A_N(net132),
    .B(net151),
    .Y(net425));
 sky130_fd_sc_hd__or3b_2 c441 (.A(net307),
    .B(net984),
    .C_N(net1001),
    .X(net426));
 sky130_fd_sc_hd__nand3b_1 c442 (.A_N(net426),
    .B(clknet_1_0__leaf_net409),
    .C(net269),
    .Y(net427));
 sky130_fd_sc_hd__clkbuf_2 c443 (.A(net908),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c444 (.A0(net133),
    .A1(net300),
    .A2(net428),
    .A3(net306),
    .S0(net426),
    .S1(net810),
    .X(net429));
 sky130_fd_sc_hd__nand3_4 c445 (.A(net307),
    .B(net428),
    .C(clknet_1_0__leaf_net427),
    .Y(net430));
 sky130_fd_sc_hd__inv_1 c446 (.A(net907),
    .Y(net431));
 sky130_fd_sc_hd__sdfsbp_2 c447 (.CLK(clknet_4_3_0_clk),
    .D(net269),
    .SCD(net428),
    .SCE(net287),
    .SET_B(net306),
    .Q(net433),
    .Q_N(net432));
 sky130_fd_sc_hd__or3b_1 c448 (.A(net425),
    .B(net290),
    .C_N(net845),
    .X(net434));
 sky130_fd_sc_hd__and3b_1 c449 (.A_N(net429),
    .B(net433),
    .C(net426),
    .X(net435));
 sky130_fd_sc_hd__and2_1 c45 (.A(net6),
    .B(net12),
    .X(net19));
 sky130_fd_sc_hd__mux4_4 c450 (.A0(net975),
    .A1(net174),
    .A2(net432),
    .A3(clknet_1_0__leaf_net427),
    .S0(net299),
    .S1(net1001),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(net412),
    .A1(net405),
    .A2(net112),
    .A3(net260),
    .S0(net432),
    .S1(net435),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net277),
    .A1(net251),
    .A2(net426),
    .A3(net412),
    .S0(net975),
    .S1(net813),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 c453 (.A(net785),
    .X(net439));
 sky130_fd_sc_hd__and2b_4 c454 (.A_N(net428),
    .B(clknet_1_0__leaf_net967),
    .X(net440));
 sky130_fd_sc_hd__or3b_1 c455 (.A(net439),
    .B(clknet_1_0__leaf_net440),
    .C_N(net1001),
    .X(net441));
 sky130_fd_sc_hd__inv_2 c456 (.A(net784),
    .Y(net442));
 sky130_fd_sc_hd__nand3_1 c457 (.A(net425),
    .B(net404),
    .C(net813),
    .Y(net443));
 sky130_fd_sc_hd__clkinv_2 c458 (.A(net829),
    .Y(net444));
 sky130_fd_sc_hd__mux4_2 c459 (.A0(net984),
    .A1(net287),
    .A2(net444),
    .A3(net260),
    .S0(clknet_1_0__leaf_net441),
    .S1(clknet_1_0__leaf_net972),
    .X(net445));
 sky130_fd_sc_hd__or2_1 c46 (.A(net938),
    .B(net930),
    .X(net20));
 sky130_fd_sc_hd__mux4_2 c460 (.A0(net443),
    .A1(net975),
    .A2(net434),
    .A3(net998),
    .S0(clknet_1_0__leaf_net409),
    .S1(net859),
    .X(net446));
 sky130_fd_sc_hd__mux4_4 c461 (.A0(net435),
    .A1(net287),
    .A2(net444),
    .A3(net432),
    .S0(clknet_1_0__leaf_net427),
    .S1(net859),
    .X(net447));
 sky130_fd_sc_hd__nor2b_1 c462 (.A(net323),
    .B_N(net309),
    .Y(net448));
 sky130_fd_sc_hd__nand2_4 c463 (.A(clknet_1_1__leaf_net427),
    .B(net325),
    .Y(net449));
 sky130_fd_sc_hd__or3b_1 c464 (.A(net442),
    .B(net46),
    .C_N(clknet_1_1__leaf_net822),
    .X(net450));
 sky130_fd_sc_hd__or4bb_1 c465 (.A(net318),
    .B(net192),
    .C_N(net231),
    .D_N(net448),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_2 c466 (.A(net816),
    .X(net452));
 sky130_fd_sc_hd__mux4_4 c467 (.A0(net323),
    .A1(clknet_1_0__leaf_net430),
    .A2(net452),
    .A3(net980),
    .S0(net934),
    .S1(clknet_1_0__leaf_net822),
    .X(net453));
 sky130_fd_sc_hd__and3b_1 c468 (.A_N(net316),
    .B(net190),
    .C(net982),
    .X(net454));
 sky130_fd_sc_hd__nand3_1 c469 (.A(net319),
    .B(net793),
    .C(net848),
    .Y(net455));
 sky130_fd_sc_hd__or2b_1 c47 (.A(net1004),
    .B_N(net19),
    .X(net21));
 sky130_fd_sc_hd__or2b_1 c470 (.A(net455),
    .B_N(net405),
    .X(net456));
 sky130_fd_sc_hd__nand2_1 c471 (.A(net456),
    .B(net167),
    .Y(net457));
 sky130_fd_sc_hd__and2_0 c472 (.A(net392),
    .B(net816),
    .X(net458));
 sky130_fd_sc_hd__nand3b_4 c473 (.A_N(clknet_1_1__leaf_net440),
    .B(net55),
    .C(clknet_1_1__leaf_net409),
    .Y(net459));
 sky130_fd_sc_hd__and3b_1 c474 (.A_N(clknet_1_1__leaf_net409),
    .B(net392),
    .C(clknet_1_0__leaf_net972),
    .X(net460));
 sky130_fd_sc_hd__nand2_4 c475 (.A(net330),
    .B(clknet_1_0__leaf_net460),
    .Y(net461));
 sky130_fd_sc_hd__mux4_2 c476 (.A0(net312),
    .A1(clknet_1_0__leaf_net461),
    .A2(clknet_1_0__leaf_net460),
    .A3(net975),
    .S0(clknet_1_1__leaf_net427),
    .S1(net308),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(clknet_1_0__leaf_net459),
    .A1(net452),
    .A2(net323),
    .A3(clknet_1_1__leaf_net460),
    .S0(net328),
    .S1(clknet_1_0__leaf_net461),
    .X(net463));
 sky130_fd_sc_hd__mux4_2 c478 (.A0(net991),
    .A1(net419),
    .A2(clknet_1_1__leaf_net460),
    .A3(net332),
    .S0(clknet_1_1__leaf_net459),
    .S1(net848),
    .X(net464));
 sky130_fd_sc_hd__mux4_4 c479 (.A0(net454),
    .A1(net457),
    .A2(clknet_1_0__leaf_net460),
    .A3(clknet_1_0__leaf_net464),
    .S0(net451),
    .S1(clknet_1_0__leaf_net461),
    .X(net465));
 sky130_fd_sc_hd__and2_1 c48 (.A(net968),
    .B(net1004),
    .X(net22));
 sky130_fd_sc_hd__nor2_2 c480 (.A(clknet_1_0__leaf_net460),
    .B(clknet_1_0__leaf_net464),
    .Y(net466));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net458),
    .A1(net457),
    .A2(clknet_1_1__leaf_net460),
    .A3(clknet_1_0__leaf_net464),
    .S0(clknet_1_0__leaf_net440),
    .S1(net865),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net430),
    .A1(clknet_1_0__leaf_net461),
    .A2(clknet_1_1__leaf_net466),
    .A3(clknet_1_0__leaf_net467),
    .S0(clknet_1_1__leaf_net460),
    .S1(net864),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net449),
    .A1(net192),
    .A2(clknet_1_0__leaf_net467),
    .A3(clknet_1_1__leaf_net409),
    .S0(clknet_1_1__leaf_net460),
    .S1(net866),
    .X(net469));
 sky130_fd_sc_hd__or4bb_1 c484 (.A(net336),
    .B(net983),
    .C_N(net1055),
    .D_N(net867),
    .X(net470));
 sky130_fd_sc_hd__or4bb_2 c485 (.A(net392),
    .B(clknet_1_0__leaf_net201),
    .C_N(net433),
    .D_N(net1003),
    .X(net471));
 sky130_fd_sc_hd__o2111ai_2 c486 (.A1(net463),
    .A2(net332),
    .B1(net987),
    .C1(net1035),
    .D1(clknet_1_0__leaf_net972),
    .Y(net472));
 sky130_fd_sc_hd__sdfbbp_1 c487 (.CLK(clknet_4_12_0_clk),
    .D(net142),
    .RESET_B(clknet_1_1__leaf_net210),
    .SCD(net1052),
    .SCE(net987),
    .SET_B(clknet_1_0__leaf_net472),
    .Q(net474),
    .Q_N(net473));
 sky130_fd_sc_hd__sdfsbp_1 c488 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net471),
    .SCD(net200),
    .SCE(net980),
    .SET_B(clknet_1_0__leaf_net967),
    .Q(net476),
    .Q_N(net475));
 sky130_fd_sc_hd__or4bb_1 c489 (.A(net192),
    .B(net419),
    .C_N(clknet_1_0__leaf_net471),
    .D_N(clknet_1_0__leaf_net472),
    .X(net477));
 sky130_fd_sc_hd__nand2_1 c49 (.A(net928),
    .B(net17),
    .Y(net23));
 sky130_fd_sc_hd__sdfstp_1 c490 (.CLK(clknet_4_14_0_clk),
    .D(net332),
    .SCD(net322),
    .SCE(net473),
    .SET_B(net866),
    .Q(net951));
 sky130_fd_sc_hd__o2111ai_2 c491 (.A1(net433),
    .A2(net356),
    .B1(clknet_1_0__leaf_net346),
    .C1(net1005),
    .D1(net475),
    .Y(net478));
 sky130_fd_sc_hd__a2111o_1 c492 (.A1(net356),
    .A2(net934),
    .B1(net433),
    .C1(net1005),
    .D1(clknet_1_1__leaf_net472),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net419),
    .A1(net476),
    .A2(net77),
    .A3(clknet_1_0__leaf_net472),
    .S0(net1005),
    .S1(net866),
    .X(net480));
 sky130_fd_sc_hd__or4bb_4 c494 (.A(clknet_1_0__leaf_net472),
    .B(net1005),
    .C_N(net332),
    .D_N(net980),
    .X(net481));
 sky130_fd_sc_hd__mux4_4 c495 (.A0(net142),
    .A1(clknet_1_1__leaf_net472),
    .A2(net328),
    .A3(net827),
    .S0(net849),
    .S1(net866),
    .X(net482));
 sky130_fd_sc_hd__sdfbbn_1 c496 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net467),
    .RESET_B(clknet_1_1__leaf_net471),
    .SCD(clknet_1_1__leaf_net472),
    .SCE(net866),
    .SET_B(net868),
    .Q(net483));
 sky130_fd_sc_hd__sdfstp_1 c497 (.CLK(clknet_4_12_0_clk),
    .D(net139),
    .SCD(net1005),
    .SCE(clknet_1_0__leaf_net472),
    .SET_B(net988),
    .Q(net484));
 sky130_fd_sc_hd__sdfstp_1 c498 (.CLK(clknet_4_6_0_clk),
    .D(net423),
    .SCD(net2),
    .SCE(net143),
    .SET_B(clknet_1_1__leaf_net472),
    .Q(net485));
 sky130_fd_sc_hd__a2111oi_0 c499 (.A1(net77),
    .A2(net980),
    .B1(net474),
    .C1(clknet_1_1__leaf_net461),
    .D1(clknet_1_1__leaf_net972),
    .Y(net486));
 sky130_fd_sc_hd__and2_1 c50 (.A(net23),
    .B(net1004),
    .X(net24));
 sky130_fd_sc_hd__sdfbbn_1 c500 (.CLK_N(clknet_4_12_0_clk),
    .D(net46),
    .RESET_B(net392),
    .SCD(clknet_1_0__leaf_net486),
    .SCE(net997),
    .SET_B(net55),
    .Q(net487));
 sky130_fd_sc_hd__sdfbbp_1 c501 (.CLK(clknet_4_12_0_clk),
    .D(net487),
    .RESET_B(clknet_1_1__leaf_net471),
    .SCD(net423),
    .SCE(net1049),
    .SET_B(net863),
    .Q(net489),
    .Q_N(net488));
 sky130_fd_sc_hd__sdfbbn_1 c502 (.CLK_N(clknet_4_12_0_clk),
    .D(net356),
    .RESET_B(clknet_1_0__leaf_net478),
    .SCD(net1000),
    .SCE(net976),
    .SET_B(net963),
    .Q(net491),
    .Q_N(net490));
 sky130_fd_sc_hd__sdfbbn_1 c503 (.CLK_N(clknet_4_12_0_clk),
    .D(net167),
    .RESET_B(net491),
    .SCD(net489),
    .SCE(net1014),
    .SET_B(clknet_1_1__leaf_net472),
    .Q(net492));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net484),
    .A1(clknet_1_1__leaf_net467),
    .A2(net490),
    .A3(net2),
    .S0(clknet_1_1__leaf_net210),
    .S1(net831),
    .X(net493));
 sky130_fd_sc_hd__mux4_4 c505 (.A0(net976),
    .A1(net483),
    .A2(net493),
    .A3(net142),
    .S0(clknet_1_1__leaf_net472),
    .S1(net488),
    .X(net494));
 sky130_fd_sc_hd__mux4_2 c509 (.A0(clknet_1_1__leaf_net201),
    .A1(net105),
    .A2(net376),
    .A3(net983),
    .S0(clknet_1_1__leaf_net841),
    .S1(clknet_1_0__leaf_net858),
    .X(net495));
 sky130_fd_sc_hd__nand2b_1 c51 (.A_N(net24),
    .B(net19),
    .Y(net25));
 sky130_fd_sc_hd__mux4_2 c510 (.A0(clknet_1_1__leaf_net241),
    .A1(net999),
    .A2(net355),
    .A3(net1005),
    .S0(net1001),
    .S1(clknet_1_1__leaf_net967),
    .X(net496));
 sky130_fd_sc_hd__mux4_2 c511 (.A0(net989),
    .A1(net983),
    .A2(net204),
    .A3(net105),
    .S0(clknet_1_1__leaf_net858),
    .S1(clknet_1_1__leaf_net967),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c512 (.A0(net355),
    .A1(net230),
    .A2(clknet_1_0__leaf_net364),
    .A3(clknet_1_1__leaf_net214),
    .S0(clknet_1_0__leaf_net841),
    .S1(net843),
    .X(net498));
 sky130_fd_sc_hd__mux4_4 c513 (.A0(net274),
    .A1(net988),
    .A2(net1005),
    .A3(clknet_1_1__leaf_net364),
    .S0(clknet_1_0__leaf_net841),
    .S1(clknet_1_1__leaf_net972),
    .X(net499));
 sky130_fd_sc_hd__mux4_4 c514 (.A0(net233),
    .A1(net204),
    .A2(clknet_1_0__leaf_net499),
    .A3(net322),
    .S0(net842),
    .S1(clknet_1_0__leaf_net858),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c515 (.A0(net230),
    .A1(net1005),
    .A2(net1000),
    .A3(net104),
    .S0(clknet_1_1__leaf_net364),
    .S1(net843),
    .X(net501));
 sky130_fd_sc_hd__mux4_4 c516 (.A0(net377),
    .A1(clknet_1_1__leaf_net499),
    .A2(clknet_1_0__leaf_net364),
    .A3(net843),
    .S0(clknet_1_1__leaf_net858),
    .S1(net871),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c517 (.A0(net498),
    .A1(net200),
    .A2(net105),
    .A3(net204),
    .S0(net980),
    .S1(net871),
    .X(net503));
 sky130_fd_sc_hd__mux4_4 c518 (.A0(net377),
    .A1(net1005),
    .A2(clknet_1_0__leaf_net499),
    .A3(clknet_1_1__leaf_net841),
    .S0(net842),
    .S1(net845),
    .X(net956));
 sky130_fd_sc_hd__mux4_4 c519 (.A0(clknet_1_1__leaf_net201),
    .A1(clknet_1_0__leaf_net501),
    .A2(clknet_1_1__leaf_net499),
    .A3(net1005),
    .S0(clknet_1_1__leaf_net364),
    .S1(net872),
    .X(net504));
 sky130_fd_sc_hd__nor2_1 c52 (.A(net20),
    .B(net23),
    .Y(net26));
 sky130_fd_sc_hd__mux4_1 c520 (.A0(net104),
    .A1(net322),
    .A2(net377),
    .A3(net355),
    .S0(clknet_1_0__leaf_net499),
    .S1(net328),
    .X(net505));
 sky130_fd_sc_hd__mux4_4 c521 (.A0(net105),
    .A1(clknet_1_1__leaf_net364),
    .A2(net104),
    .A3(net867),
    .S0(net872),
    .S1(net873),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c522 (.A0(net287),
    .A1(net350),
    .A2(net230),
    .A3(clknet_1_1__leaf_net858),
    .S0(net871),
    .S1(net873),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(net322),
    .A1(net274),
    .A2(net376),
    .A3(net1000),
    .S0(net867),
    .S1(net1046),
    .X(net508));
 sky130_fd_sc_hd__mux4_4 c524 (.A0(clknet_1_1__leaf_net364),
    .A1(clknet_1_0__leaf_net502),
    .A2(clknet_1_1__leaf_net499),
    .A3(clknet_1_0__leaf_net501),
    .S0(net872),
    .S1(net873),
    .X(net509));
 sky130_fd_sc_hd__mux4_4 c525 (.A0(clknet_1_1__leaf_net502),
    .A1(net1000),
    .A2(net355),
    .A3(net807),
    .S0(net870),
    .S1(net873),
    .X(net510));
 sky130_fd_sc_hd__mux4_2 c526 (.A0(net504),
    .A1(clknet_1_1__leaf_net501),
    .A2(net981),
    .A3(net867),
    .S0(net873),
    .S1(clknet_1_0__leaf_net875),
    .X(net511));
 sky130_fd_sc_hd__mux4_2 c527 (.A0(net1013),
    .A1(clknet_1_1__leaf_net364),
    .A2(net826),
    .A3(net872),
    .S0(net874),
    .S1(clknet_1_1__leaf_net875),
    .X(net965));
 sky130_fd_sc_hd__nand2_4 c528 (.A(net923),
    .B(net112),
    .Y(net512));
 sky130_fd_sc_hd__inv_4 c529 (.A(net742),
    .Y(net513));
 sky130_fd_sc_hd__or2b_1 c53 (.A(net26),
    .B_N(net20),
    .X(net27));
 sky130_fd_sc_hd__nor2_1 c530 (.A(net512),
    .B(net401),
    .Y(net514));
 sky130_fd_sc_hd__buf_1 c531 (.A(net742),
    .X(net515));
 sky130_fd_sc_hd__and2b_1 c532 (.A_N(net926),
    .B(net388),
    .X(net516));
 sky130_fd_sc_hd__nand2b_2 c533 (.A_N(net516),
    .B(net381),
    .Y(net517));
 sky130_fd_sc_hd__or2b_1 c534 (.A(net1062),
    .B_N(net825),
    .X(net518));
 sky130_fd_sc_hd__nand2b_4 c535 (.A_N(net260),
    .B(net515),
    .Y(net519));
 sky130_fd_sc_hd__inv_4 c536 (.A(net769),
    .Y(net520));
 sky130_fd_sc_hd__buf_1 c537 (.A(net774),
    .X(net521));
 sky130_fd_sc_hd__and2b_2 c538 (.A_N(net397),
    .B(net520),
    .X(net522));
 sky130_fd_sc_hd__inv_4 c539 (.A(net774),
    .Y(net523));
 sky130_fd_sc_hd__nand2_1 c54 (.A(net27),
    .B(net938),
    .Y(net28));
 sky130_fd_sc_hd__nand2b_1 c540 (.A_N(net522),
    .B(net516),
    .Y(net524));
 sky130_fd_sc_hd__sedfxbp_2 c541 (.CLK(clknet_4_1_0_clk),
    .D(net264),
    .DE(net514),
    .SCD(net518),
    .SCE(net517),
    .Q(net526),
    .Q_N(net525));
 sky130_fd_sc_hd__and2_2 c542 (.A(net524),
    .B(net381),
    .X(net527));
 sky130_fd_sc_hd__sedfxbp_1 c543 (.CLK(clknet_4_1_0_clk),
    .D(net1062),
    .DE(net383),
    .SCD(net525),
    .SCE(net246),
    .Q(net529),
    .Q_N(net528));
 sky130_fd_sc_hd__a2111o_1 c544 (.A1(net517),
    .A2(net384),
    .B1(net527),
    .C1(net512),
    .D1(net514),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net520),
    .A1(net527),
    .A2(net517),
    .A3(net381),
    .S0(net384),
    .S1(net825),
    .X(net531));
 sky130_fd_sc_hd__mux4_2 c546 (.A0(net522),
    .A1(net528),
    .A2(net524),
    .A3(net525),
    .S0(net254),
    .S1(clknet_1_0__leaf_net876),
    .X(net532));
 sky130_fd_sc_hd__or4bb_4 c547 (.A(net516),
    .B(clknet_1_0__leaf_net532),
    .C_N(net805),
    .D_N(clknet_1_0__leaf_net876),
    .X(net533));
 sky130_fd_sc_hd__or4bb_4 c548 (.A(clknet_1_0__leaf_net532),
    .B(clknet_1_0__leaf_net533),
    .C_N(net519),
    .D_N(clknet_1_1__leaf_net876),
    .X(net534));
 sky130_fd_sc_hd__mux4_4 c549 (.A0(net246),
    .A1(clknet_1_0__leaf_net534),
    .A2(net517),
    .A3(clknet_1_0__leaf_net533),
    .S0(net522),
    .S1(clknet_1_1__leaf_net876),
    .X(net535));
 sky130_fd_sc_hd__nor2_2 c55 (.A(net18),
    .B(net19),
    .Y(net29));
 sky130_fd_sc_hd__inv_2 c550 (.A(net817),
    .Y(net536));
 sky130_fd_sc_hd__or3b_4 c551 (.A(net941),
    .B(net936),
    .C_N(net846),
    .X(net537));
 sky130_fd_sc_hd__buf_6 c552 (.A(net817),
    .X(net538));
 sky130_fd_sc_hd__nand3_2 c553 (.A(net391),
    .B(net537),
    .C(net538),
    .Y(net539));
 sky130_fd_sc_hd__or3_4 c554 (.A(net529),
    .B(clknet_1_1__leaf_net533),
    .C(net268),
    .X(net540));
 sky130_fd_sc_hd__and2b_1 c555 (.A_N(net4),
    .B(net519),
    .X(net541));
 sky130_fd_sc_hd__and2_2 c556 (.A(net413),
    .B(net541),
    .X(net542));
 sky130_fd_sc_hd__and2_1 c557 (.A(net384),
    .B(net4),
    .X(net543));
 sky130_fd_sc_hd__nor2b_1 c558 (.A(net539),
    .B_N(net523),
    .Y(net544));
 sky130_fd_sc_hd__nand3b_1 c559 (.A_N(net272),
    .B(net413),
    .C(net121),
    .Y(net545));
 sky130_fd_sc_hd__nor2b_1 c56 (.A(net25),
    .B_N(net20),
    .Y(net30));
 sky130_fd_sc_hd__and3_1 c560 (.A(net421),
    .B(net413),
    .C(net545),
    .X(net546));
 sky130_fd_sc_hd__nor2b_2 c561 (.A(net518),
    .B_N(net121),
    .Y(net547));
 sky130_fd_sc_hd__or3b_4 c562 (.A(clknet_1_1__leaf_net533),
    .B(net1032),
    .C_N(net272),
    .X(net548));
 sky130_fd_sc_hd__or4bb_2 c563 (.A(net415),
    .B(clknet_1_0__leaf_net548),
    .C_N(clknet_1_1__leaf_net540),
    .D_N(net542),
    .X(net549));
 sky130_fd_sc_hd__and3b_1 c564 (.A_N(net514),
    .B(net547),
    .C(net538),
    .X(net550));
 sky130_fd_sc_hd__nand3b_4 c565 (.A_N(net541),
    .B(net2),
    .C(net539),
    .Y(net551));
 sky130_fd_sc_hd__inv_1 c566 (.A(net922),
    .Y(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 c567 (.A(net817),
    .X(net553));
 sky130_fd_sc_hd__mux4_2 c568 (.A0(clknet_1_1__leaf_net420),
    .A1(net542),
    .A2(net551),
    .A3(clknet_1_0__leaf_net548),
    .S0(net254),
    .S1(net260),
    .X(net554));
 sky130_fd_sc_hd__buf_1 c569 (.A(net817),
    .X(net555));
 sky130_fd_sc_hd__nor2b_1 c57 (.A(net5),
    .B_N(net24),
    .Y(net31));
 sky130_fd_sc_hd__mux4_2 c570 (.A0(net545),
    .A1(clknet_1_0__leaf_net540),
    .A2(net551),
    .A3(net538),
    .S0(net251),
    .S1(clknet_1_0__leaf_net533),
    .X(net556));
 sky130_fd_sc_hd__mux4_2 c571 (.A0(net553),
    .A1(net551),
    .A2(net537),
    .A3(net143),
    .S0(clknet_1_0__leaf_net548),
    .S1(net545),
    .X(net557));
 sky130_fd_sc_hd__nand2_1 c572 (.A(net260),
    .B(net300),
    .Y(net558));
 sky130_fd_sc_hd__or4bb_1 c573 (.A(net251),
    .B(net975),
    .C_N(net558),
    .D_N(net860),
    .X(net559));
 sky130_fd_sc_hd__or4bb_1 c574 (.A(net434),
    .B(net260),
    .C_N(net405),
    .D_N(net941),
    .X(net560));
 sky130_fd_sc_hd__and2_0 c575 (.A(net155),
    .B(net308),
    .X(net561));
 sky130_fd_sc_hd__nand3b_2 c576 (.A_N(net173),
    .B(net847),
    .C(clknet_1_0__leaf_net967),
    .Y(net562));
 sky130_fd_sc_hd__sedfxtp_4 c577 (.CLK(clknet_4_1_0_clk),
    .D(net558),
    .DE(net403),
    .SCD(net251),
    .SCE(net975),
    .Q(net563));
 sky130_fd_sc_hd__dlymetal6s2s_1 c578 (.A(net909),
    .X(net564));
 sky130_fd_sc_hd__mux4_2 c579 (.A0(net174),
    .A1(net990),
    .A2(net527),
    .A3(net563),
    .S0(net299),
    .S1(clknet_1_0__leaf_net562),
    .X(net565));
 sky130_fd_sc_hd__nand2_1 c58 (.A(net6),
    .B(net25),
    .Y(net32));
 sky130_fd_sc_hd__sedfxtp_2 c580 (.CLK(clknet_4_1_0_clk),
    .D(net527),
    .DE(net444),
    .SCD(net975),
    .SCE(net563),
    .Q(net566));
 sky130_fd_sc_hd__or4bb_1 c581 (.A(net112),
    .B(net444),
    .C_N(net512),
    .D_N(net404),
    .X(net567));
 sky130_fd_sc_hd__and3_1 c582 (.A(net251),
    .B(net112),
    .C(net566),
    .X(net568));
 sky130_fd_sc_hd__mux4_4 c583 (.A0(net567),
    .A1(net561),
    .A2(net566),
    .A3(clknet_1_0__leaf_net441),
    .S0(clknet_1_0__leaf_net562),
    .S1(net1000),
    .X(net569));
 sky130_fd_sc_hd__or4bb_1 c584 (.A(net2),
    .B(net566),
    .C_N(net564),
    .D_N(net877),
    .X(net570));
 sky130_fd_sc_hd__a2111o_1 c585 (.A1(net546),
    .A2(net563),
    .B1(net112),
    .C1(net941),
    .D1(net878),
    .X(net571));
 sky130_fd_sc_hd__and2b_1 c586 (.A_N(net570),
    .B(net563),
    .X(net572));
 sky130_fd_sc_hd__o2111a_1 c587 (.A1(net571),
    .A2(net564),
    .B1(net860),
    .C1(net861),
    .D1(net878),
    .X(net573));
 sky130_fd_sc_hd__or4bb_1 c588 (.A(net566),
    .B(net563),
    .C_N(clknet_1_0__leaf_net562),
    .D_N(net546),
    .X(net574));
 sky130_fd_sc_hd__or4bb_1 c589 (.A(net431),
    .B(net112),
    .C_N(net260),
    .D_N(net877),
    .X(net950));
 sky130_fd_sc_hd__mux4_1 c59 (.A0(net937),
    .A1(net14),
    .A2(net32),
    .A3(net31),
    .S0(net924),
    .S1(net1004),
    .X(net33));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net573),
    .A1(net566),
    .A2(net563),
    .A3(net444),
    .S0(net997),
    .S1(net878),
    .X(net575));
 sky130_fd_sc_hd__mux4_2 c591 (.A0(net551),
    .A1(clknet_1_0__leaf_net574),
    .A2(net547),
    .A3(net564),
    .S0(net877),
    .S1(net879),
    .X(net576));
 sky130_fd_sc_hd__mux4_2 c592 (.A0(clknet_1_0__leaf_net441),
    .A1(net431),
    .A2(net564),
    .A3(clknet_1_0__leaf_net574),
    .S0(net847),
    .S1(net862),
    .X(net577));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net560),
    .A1(net142),
    .A2(net147),
    .A3(net173),
    .S0(clknet_1_0__leaf_net574),
    .S1(net879),
    .X(net578));
 sky130_fd_sc_hd__or4bb_4 c594 (.A(net526),
    .B(clknet_1_0__leaf_net557),
    .C_N(net542),
    .D_N(net299),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net190),
    .A1(net551),
    .A2(net448),
    .A3(clknet_1_0__leaf_net464),
    .S0(net299),
    .S1(clknet_1_0__leaf_net441),
    .X(net580));
 sky130_fd_sc_hd__or4bb_1 c596 (.A(net450),
    .B(clknet_1_0__leaf_net464),
    .C_N(net564),
    .D_N(net547),
    .X(net581));
 sky130_fd_sc_hd__and3b_1 c597 (.A_N(net405),
    .B(net980),
    .C(net1044),
    .X(net582));
 sky130_fd_sc_hd__o2111a_2 c598 (.A1(net568),
    .A2(clknet_1_0__leaf_net466),
    .B1(clknet_1_0__leaf_net441),
    .C1(clknet_1_1__leaf_net579),
    .D1(net867),
    .X(net583));
 sky130_fd_sc_hd__or4bb_2 c599 (.A(net300),
    .B(net1035),
    .C_N(clknet_1_0__leaf_net441),
    .D_N(net999),
    .X(net584));
 sky130_fd_sc_hd__and2b_1 c60 (.A_N(net30),
    .B(net25),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 c600 (.A(net744),
    .X(net585));
 sky130_fd_sc_hd__or4bb_1 c601 (.A(net527),
    .B(clknet_1_1__leaf_net441),
    .C_N(clknet_1_0__leaf_net821),
    .D_N(net877),
    .X(net586));
 sky130_fd_sc_hd__sedfxtp_4 c602 (.CLK(clknet_4_6_0_clk),
    .D(net547),
    .DE(clknet_1_0__leaf_net466),
    .SCD(clknet_1_0__leaf_net461),
    .SCE(clknet_1_1__leaf_net583),
    .Q(net587));
 sky130_fd_sc_hd__buf_6 c603 (.A(net743),
    .X(net588));
 sky130_fd_sc_hd__sdfbbp_1 c604 (.CLK(clknet_4_6_0_clk),
    .D(net588),
    .RESET_B(clknet_1_1__leaf_net557),
    .SCD(clknet_1_0__leaf_net583),
    .SCE(net547),
    .SET_B(net878),
    .Q(net590),
    .Q_N(net589));
 sky130_fd_sc_hd__sdfbbn_2 c605 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net579),
    .RESET_B(clknet_1_0__leaf_net584),
    .SCD(clknet_1_0__leaf_net557),
    .SCE(clknet_1_0__leaf_net583),
    .SET_B(net1040),
    .Q(net949),
    .Q_N(net591));
 sky130_fd_sc_hd__o2111a_1 c606 (.A1(net448),
    .A2(net526),
    .B1(clknet_1_1__leaf_net584),
    .C1(net300),
    .D1(net998),
    .X(net592));
 sky130_fd_sc_hd__or4bb_4 c607 (.A(net564),
    .B(clknet_1_0__leaf_net581),
    .C_N(net591),
    .D_N(net999),
    .X(net957));
 sky130_fd_sc_hd__nand3b_4 c608 (.A_N(clknet_1_1__leaf_net466),
    .B(net587),
    .C(net325),
    .Y(net593));
 sky130_fd_sc_hd__mux4_4 c609 (.A0(net592),
    .A1(net949),
    .A2(net526),
    .A3(net980),
    .S0(net537),
    .S1(clknet_1_0__leaf_net593),
    .X(net594));
 sky130_fd_sc_hd__nor2b_1 c61 (.A(net941),
    .B_N(net6),
    .Y(net35));
 sky130_fd_sc_hd__mux4_4 c610 (.A0(net585),
    .A1(clknet_1_1__leaf_net593),
    .A2(net589),
    .A3(net591),
    .S0(net319),
    .S1(net881),
    .X(net595));
 sky130_fd_sc_hd__mux4_4 c611 (.A0(net551),
    .A1(net590),
    .A2(net55),
    .A3(clknet_1_0__leaf_net580),
    .S0(clknet_1_1__leaf_net593),
    .S1(net802),
    .X(net596));
 sky130_fd_sc_hd__mux4_4 c612 (.A0(net924),
    .A1(net527),
    .A2(net588),
    .A3(clknet_1_1__leaf_net593),
    .S0(net200),
    .S1(net883),
    .X(net597));
 sky130_fd_sc_hd__sdfrbp_1 c613 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_0__leaf_net593),
    .RESET_B(net582),
    .SCD(net319),
    .SCE(net882),
    .Q(net599),
    .Q_N(net598));
 sky130_fd_sc_hd__mux4_2 c614 (.A0(net572),
    .A1(clknet_1_0__leaf_net593),
    .A2(net582),
    .A3(clknet_1_0__leaf_net461),
    .S0(clknet_1_1__leaf_net581),
    .S1(net883),
    .X(net600));
 sky130_fd_sc_hd__o2111a_1 c615 (.A1(net200),
    .A2(net588),
    .B1(net802),
    .C1(net1041),
    .D1(net1051),
    .X(net601));
 sky130_fd_sc_hd__sdfbbn_1 c616 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net210),
    .RESET_B(clknet_1_1__leaf_net578),
    .SCD(net489),
    .SCE(net934),
    .SET_B(net1041),
    .Q(net960),
    .Q_N(net602));
 sky130_fd_sc_hd__o2111a_4 c617 (.A1(net489),
    .A2(net143),
    .B1(clknet_1_0__leaf_net578),
    .C1(net602),
    .D1(net204),
    .X(net603));
 sky130_fd_sc_hd__mux4_4 c618 (.A0(clknet_1_1__leaf_net580),
    .A1(net997),
    .A2(net987),
    .A3(net1012),
    .S0(net328),
    .S1(clknet_1_1__leaf_net972),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net55),
    .A1(net537),
    .A2(clknet_1_0__leaf_net580),
    .A3(net981),
    .S0(net1003),
    .S1(net952),
    .X(net605));
 sky130_fd_sc_hd__or2b_1 c62 (.A(net33),
    .B_N(net21),
    .X(net36));
 sky130_fd_sc_hd__a2111o_1 c620 (.A1(net519),
    .A2(net143),
    .B1(net473),
    .C1(net1003),
    .D1(net961),
    .X(net969));
 sky130_fd_sc_hd__o2111ai_4 c621 (.A1(clknet_1_1__leaf_net346),
    .A2(net519),
    .B1(net150),
    .C1(net882),
    .D1(net961),
    .Y(net606));
 sky130_fd_sc_hd__sdfbbp_1 c622 (.CLK(clknet_4_6_0_clk),
    .D(net576),
    .RESET_B(net527),
    .SCD(net1000),
    .SCE(net934),
    .SET_B(net1048),
    .Q(net608),
    .Q_N(net607));
 sky130_fd_sc_hd__sdfbbn_1 c623 (.CLK_N(clknet_4_13_0_clk),
    .D(net537),
    .RESET_B(net1058),
    .SCD(net587),
    .SCE(net975),
    .SET_B(net961),
    .Q(net610),
    .Q_N(net609));
 sky130_fd_sc_hd__a2111o_4 c624 (.A1(net492),
    .A2(net608),
    .B1(clknet_1_1__leaf_net461),
    .C1(net928),
    .D1(net812),
    .X(net611));
 sky130_fd_sc_hd__a2111o_1 c625 (.A1(net590),
    .A2(clknet_1_0__leaf_net611),
    .B1(clknet_1_1__leaf_net210),
    .C1(net607),
    .D1(net961),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net474),
    .A1(clknet_1_1__leaf_net461),
    .A2(clknet_1_0__leaf_net611),
    .A3(net960),
    .S0(net609),
    .S1(clknet_1_0__leaf_net346),
    .X(net613));
 sky130_fd_sc_hd__o2111ai_2 c627 (.A1(net966),
    .A2(clknet_1_1__leaf_net611),
    .B1(clknet_1_1__leaf_net461),
    .C1(clknet_1_1__leaf_net821),
    .D1(clknet_1_1__leaf_net967),
    .Y(net614));
 sky130_fd_sc_hd__sdfbbn_1 c628 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net613),
    .RESET_B(net601),
    .SCD(net591),
    .SCE(clknet_1_0__leaf_net957),
    .SET_B(net527),
    .Q(net616),
    .Q_N(net615));
 sky130_fd_sc_hd__o2111ai_2 c629 (.A1(net606),
    .A2(net616),
    .B1(net966),
    .C1(clknet_1_0__leaf_net611),
    .D1(net607),
    .Y(net617));
 sky130_fd_sc_hd__mux4_1 c63 (.A0(net34),
    .A1(net6),
    .A2(net24),
    .A3(net29),
    .S0(net30),
    .S1(net25),
    .X(net37));
 sky130_fd_sc_hd__sdfbbp_1 c630 (.CLK(clknet_4_6_0_clk),
    .D(net1043),
    .RESET_B(net612),
    .SCD(net1059),
    .SCE(net537),
    .SET_B(net849),
    .Q(net618));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(clknet_1_1__leaf_net478),
    .A1(net618),
    .A2(net610),
    .A3(net608),
    .S0(net1036),
    .S1(net881),
    .X(net619));
 sky130_fd_sc_hd__o2111a_2 c632 (.A1(net587),
    .A2(net616),
    .B1(net1011),
    .C1(clknet_1_1__leaf_net461),
    .D1(net607),
    .X(net620));
 sky130_fd_sc_hd__a2111oi_2 c633 (.A1(net620),
    .A2(clknet_1_1__leaf_net611),
    .B1(net615),
    .C1(net812),
    .D1(clknet_1_1__leaf_net972),
    .Y(net621));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net577),
    .A1(net610),
    .A2(clknet_1_0__leaf_net621),
    .A3(clknet_1_1__leaf_net611),
    .S0(net987),
    .S1(net1001),
    .X(net622));
 sky130_fd_sc_hd__o2111a_2 c635 (.A1(net608),
    .A2(net614),
    .B1(clknet_1_1__leaf_net613),
    .C1(clknet_1_1__leaf_net611),
    .D1(net867),
    .X(net623));
 sky130_fd_sc_hd__mux4_2 c636 (.A0(net623),
    .A1(net608),
    .A2(clknet_1_1__leaf_net461),
    .A3(net971),
    .S0(net961),
    .S1(net884),
    .X(net624));
 sky130_fd_sc_hd__a2111oi_4 c637 (.A1(net624),
    .A2(clknet_1_1__leaf_net621),
    .B1(net1010),
    .C1(net987),
    .D1(net609),
    .Y(net625));
 sky130_fd_sc_hd__or2_1 c64 (.A(net30),
    .B(net28),
    .X(net38));
 sky130_fd_sc_hd__and2_1 c65 (.A(net933),
    .B(net928),
    .X(net39));
 sky130_fd_sc_hd__and2b_1 c66 (.A_N(net21),
    .B(net18),
    .X(net40));
 sky130_fd_sc_hd__nor2_1 c660 (.A(net925),
    .B(net401),
    .Y(net626));
 sky130_fd_sc_hd__and2b_1 c661 (.A_N(net526),
    .B(net389),
    .X(net627));
 sky130_fd_sc_hd__nor2b_1 c662 (.A(net521),
    .B_N(net522),
    .Y(net628));
 sky130_fd_sc_hd__nor2b_1 c663 (.A(net936),
    .B_N(clknet_1_0__leaf_net534),
    .Y(net629));
 sky130_fd_sc_hd__or2b_1 c664 (.A(net381),
    .B_N(net994),
    .X(net630));
 sky130_fd_sc_hd__and2b_1 c665 (.A_N(net513),
    .B(net519),
    .X(net631));
 sky130_fd_sc_hd__or2b_1 c666 (.A(net994),
    .B_N(net513),
    .X(net632));
 sky130_fd_sc_hd__nor2_4 c667 (.A(net931),
    .B(net994),
    .Y(net633));
 sky130_fd_sc_hd__inv_4 c668 (.A(net820),
    .Y(net634));
 sky130_fd_sc_hd__and2b_1 c669 (.A_N(net632),
    .B(net512),
    .X(net635));
 sky130_fd_sc_hd__or2_1 c67 (.A(net933),
    .B(net982),
    .X(net41));
 sky130_fd_sc_hd__nor2b_2 c670 (.A(net634),
    .B_N(net521),
    .Y(net636));
 sky130_fd_sc_hd__nor2b_1 c671 (.A(net636),
    .B_N(net525),
    .Y(net637));
 sky130_fd_sc_hd__nor2b_2 c672 (.A(net631),
    .B_N(net636),
    .Y(net638));
 sky130_fd_sc_hd__and3_2 c673 (.A(net638),
    .B(net521),
    .C(clknet_1_0__leaf_net629),
    .X(net639));
 sky130_fd_sc_hd__nand2_2 c674 (.A(clknet_1_1__leaf_net629),
    .B(net638),
    .Y(net640));
 sky130_fd_sc_hd__or3_2 c675 (.A(net388),
    .B(net638),
    .C(clknet_1_0__leaf_net639),
    .X(net641));
 sky130_fd_sc_hd__or3_4 c676 (.A(net627),
    .B(net401),
    .C(net638),
    .X(net642));
 sky130_fd_sc_hd__nand3_4 c677 (.A(net642),
    .B(net633),
    .C(net638),
    .Y(net643));
 sky130_fd_sc_hd__clkbuf_1 c678 (.A(net820),
    .X(net644));
 sky130_fd_sc_hd__and3_4 c679 (.A(clknet_1_1__leaf_net534),
    .B(net642),
    .C(net633),
    .X(net645));
 sky130_fd_sc_hd__nor2b_1 c68 (.A(net31),
    .B_N(net40),
    .Y(net42));
 sky130_fd_sc_hd__a2111o_4 c680 (.A1(net644),
    .A2(clknet_1_0__leaf_net641),
    .B1(net642),
    .C1(net637),
    .D1(net643),
    .X(net646));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net634),
    .A1(net636),
    .A2(net642),
    .A3(net633),
    .S0(net630),
    .S1(net805),
    .X(net647));
 sky130_fd_sc_hd__o2111a_2 c682 (.A1(net389),
    .A2(net404),
    .B1(clknet_1_1__leaf_net645),
    .C1(net635),
    .D1(net847),
    .X(net648));
 sky130_fd_sc_hd__nor3b_2 c683 (.A(clknet_1_1__leaf_net556),
    .B(net555),
    .C_N(net538),
    .Y(net649));
 sky130_fd_sc_hd__sdfrbp_1 c684 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net645),
    .RESET_B(net1054),
    .SCD(net522),
    .SCE(net1007),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__or3_2 c685 (.A(net523),
    .B(net651),
    .C(net403),
    .X(net652));
 sky130_fd_sc_hd__sdfrtn_1 c686 (.CLK_N(clknet_4_4_0_clk),
    .D(net536),
    .RESET_B(clknet_1_1__leaf_net641),
    .SCD(net401),
    .SCE(net801),
    .Q(net653));
 sky130_fd_sc_hd__nand3b_4 c687 (.A_N(net636),
    .B(net150),
    .C(net650),
    .Y(net654));
 sky130_fd_sc_hd__o2111a_2 c688 (.A1(net401),
    .A2(clknet_1_1__leaf_net548),
    .B1(clknet_1_0__leaf_net556),
    .C1(net522),
    .D1(net653),
    .X(net655));
 sky130_fd_sc_hd__inv_4 c689 (.A(net740),
    .Y(net656));
 sky130_fd_sc_hd__and2_1 c69 (.A(net40),
    .B(net939),
    .X(net43));
 sky130_fd_sc_hd__and3b_2 c690 (.A_N(net940),
    .B(clknet_1_0__leaf_net655),
    .C(net654),
    .X(net657));
 sky130_fd_sc_hd__nor3b_2 c691 (.A(clknet_1_1__leaf_net649),
    .B(net522),
    .C_N(net820),
    .Y(net658));
 sky130_fd_sc_hd__clkbuf_2 c692 (.A(net739),
    .X(net659));
 sky130_fd_sc_hd__buf_4 c693 (.A(clknet_1_1__leaf_net912),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__nor3_4 c695 (.A(net651),
    .B(net660),
    .C(net656),
    .Y(net662));
 sky130_fd_sc_hd__a2111oi_0 c696 (.A1(clknet_1_1__leaf_net662),
    .A2(net656),
    .B1(net633),
    .C1(net653),
    .D1(net637),
    .Y(net663));
 sky130_fd_sc_hd__o2111ai_4 c697 (.A1(clknet_1_1__leaf_net533),
    .A2(clknet_1_0__leaf_net662),
    .B1(net654),
    .C1(net403),
    .D1(net404),
    .Y(net664));
 sky130_fd_sc_hd__a2111o_2 c698 (.A1(net654),
    .A2(clknet_1_0__leaf_net662),
    .B1(net650),
    .C1(clknet_1_1__leaf_net548),
    .D1(net801),
    .X(net665));
 sky130_fd_sc_hd__mux4_2 c699 (.A0(net552),
    .A1(clknet_1_1__leaf_net655),
    .A2(clknet_1_0__leaf_net649),
    .A3(clknet_1_0__leaf_net662),
    .S0(clknet_1_1__leaf_net548),
    .S1(net653),
    .X(net666));
 sky130_fd_sc_hd__nor2b_1 c70 (.A(net36),
    .B_N(net29),
    .Y(net44));
 sky130_fd_sc_hd__mux4_2 c700 (.A0(net628),
    .A1(net663),
    .A2(clknet_1_0__leaf_net664),
    .A3(clknet_1_1__leaf_net662),
    .S0(net404),
    .S1(net538),
    .X(net667));
 sky130_fd_sc_hd__sdfbbn_1 c701 (.CLK_N(clknet_4_5_0_clk),
    .D(net538),
    .RESET_B(net1033),
    .SCD(clknet_1_0__leaf_net664),
    .SCE(clknet_1_0__leaf_net665),
    .SET_B(net800),
    .Q(net669),
    .Q_N(net668));
 sky130_fd_sc_hd__mux4_2 c702 (.A0(net658),
    .A1(net637),
    .A2(net643),
    .A3(net653),
    .S0(net636),
    .S1(net885),
    .X(net670));
 sky130_fd_sc_hd__sdfbbn_1 c703 (.CLK_N(clknet_4_5_0_clk),
    .D(clknet_1_1__leaf_net657),
    .RESET_B(net1042),
    .SCD(net1007),
    .SCE(clknet_1_1__leaf_net662),
    .SET_B(net800),
    .Q(net672),
    .Q_N(net671));
 sky130_fd_sc_hd__sdfrtp_1 c704 (.CLK(clknet_4_4_0_clk),
    .D(net404),
    .RESET_B(clknet_1_0__leaf_net666),
    .SCD(net519),
    .SCE(clknet_1_0__leaf_net554),
    .Q(net673));
 sky130_fd_sc_hd__nand3b_2 c705 (.A_N(net403),
    .B(clknet_1_0__leaf_net562),
    .C(net846),
    .Y(net674));
 sky130_fd_sc_hd__and3_1 c706 (.A(net635),
    .B(net308),
    .C(net880),
    .X(net675));
 sky130_fd_sc_hd__nand3_2 c707 (.A(net673),
    .B(net659),
    .C(net880),
    .Y(net676));
 sky130_fd_sc_hd__or4bb_1 c708 (.A(net640),
    .B(net403),
    .C_N(net404),
    .D_N(net847),
    .X(net677));
 sky130_fd_sc_hd__a2111o_4 c709 (.A1(net659),
    .A2(clknet_1_1__leaf_net554),
    .B1(net147),
    .C1(net519),
    .D1(net668),
    .X(net678));
 sky130_fd_sc_hd__inv_6 c71 (.A(net751),
    .Y(net45));
 sky130_fd_sc_hd__nor3_1 c710 (.A(net444),
    .B(clknet_1_0__leaf_net562),
    .C(clknet_1_1__leaf_net574),
    .Y(net679));
 sky130_fd_sc_hd__o2111ai_4 c711 (.A1(net659),
    .A2(clknet_1_0__leaf_net664),
    .B1(net984),
    .C1(clknet_1_0__leaf_net562),
    .D1(net968),
    .Y(net680));
 sky130_fd_sc_hd__a2111o_4 c712 (.A1(clknet_1_1__leaf_net574),
    .A2(net1007),
    .B1(clknet_1_0__leaf_net678),
    .C1(net308),
    .D1(net928),
    .X(net681));
 sky130_fd_sc_hd__and3_1 c713 (.A(net654),
    .B(net147),
    .C(net879),
    .X(net682));
 sky130_fd_sc_hd__a2111oi_4 c714 (.A1(clknet_1_1__leaf_net548),
    .A2(net676),
    .B1(net654),
    .C1(net643),
    .D1(net525),
    .Y(net683));
 sky130_fd_sc_hd__sdfbbp_1 c715 (.CLK(clknet_4_4_0_clk),
    .D(net924),
    .RESET_B(clknet_1_0__leaf_net674),
    .SCD(clknet_1_0__leaf_net678),
    .SCE(net847),
    .SET_B(net880),
    .Q(net685),
    .Q_N(net684));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net673),
    .A1(net404),
    .A2(net669),
    .A3(clknet_1_1__leaf_net664),
    .S0(net563),
    .S1(net444),
    .X(net686));
 sky130_fd_sc_hd__buf_16 c717 (.A(net909),
    .X(net687));
 sky130_fd_sc_hd__o2111ai_1 c718 (.A1(net626),
    .A2(net682),
    .B1(net519),
    .C1(net846),
    .D1(net889),
    .Y(net688));
 sky130_fd_sc_hd__sdfbbn_2 c719 (.CLK_N(clknet_4_4_0_clk),
    .D(clknet_1_1__leaf_net666),
    .RESET_B(net404),
    .SCD(net684),
    .SCE(net830),
    .SET_B(net889),
    .Q(net690),
    .Q_N(net689));
 sky130_fd_sc_hd__clkbuf_2 c72 (.A(net751),
    .X(net46));
 sky130_fd_sc_hd__nor3_1 c720 (.A(net675),
    .B(net984),
    .C(net889),
    .Y(net691));
 sky130_fd_sc_hd__sdfbbn_2 c721 (.CLK_N(clknet_4_5_0_clk),
    .D(net147),
    .RESET_B(clknet_1_1__leaf_net574),
    .SCD(clknet_1_1__leaf_net678),
    .SCE(net643),
    .SET_B(net563),
    .Q(net693),
    .Q_N(net692));
 sky130_fd_sc_hd__sdfbbp_1 c722 (.CLK(clknet_4_5_0_clk),
    .D(net688),
    .RESET_B(clknet_1_1__leaf_net678),
    .SCD(net689),
    .SCE(net685),
    .SET_B(net692),
    .Q(net695),
    .Q_N(net694));
 sky130_fd_sc_hd__a2111o_4 c723 (.A1(net669),
    .A2(net695),
    .B1(net687),
    .C1(net889),
    .D1(clknet_1_1__leaf_net678),
    .X(net696));
 sky130_fd_sc_hd__o2111ai_4 c724 (.A1(net681),
    .A2(net691),
    .B1(net690),
    .C1(net692),
    .D1(clknet_1_1__leaf_net664),
    .Y(net697));
 sky130_fd_sc_hd__sdfbbn_1 c725 (.CLK_N(clknet_4_5_0_clk),
    .D(net643),
    .RESET_B(net1047),
    .SCD(clknet_1_0__leaf_net696),
    .SCE(net830),
    .SET_B(net889),
    .Q(net699),
    .Q_N(net698));
 sky130_fd_sc_hd__mux4_2 c726 (.A0(net542),
    .A1(net693),
    .A2(clknet_1_0__leaf_net674),
    .A3(net694),
    .S0(net689),
    .S1(net319),
    .X(net700));
 sky130_fd_sc_hd__a2111oi_4 c727 (.A1(clknet_1_1__leaf_net441),
    .A2(net997),
    .B1(clknet_1_0__leaf_net679),
    .C1(net598),
    .D1(net684),
    .Y(net701));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net695),
    .A1(net693),
    .A2(net1007),
    .A3(net815),
    .S0(net885),
    .S1(net887),
    .X(net702));
 sky130_fd_sc_hd__sdfbbn_1 c729 (.CLK_N(clknet_4_5_0_clk),
    .D(net633),
    .RESET_B(net309),
    .SCD(clknet_1_0__leaf_net674),
    .SCE(net692),
    .SET_B(clknet_1_1__leaf_net562),
    .Q(net703));
 sky130_fd_sc_hd__and2_1 c73 (.A(net45),
    .B(net28),
    .X(net47));
 sky130_fd_sc_hd__mux4_4 c730 (.A0(clknet_1_1__leaf_net562),
    .A1(net542),
    .A2(net687),
    .A3(net671),
    .S0(net849),
    .S1(net865),
    .X(net704));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net599),
    .A1(net633),
    .A2(net690),
    .A3(clknet_1_1__leaf_net696),
    .S0(clknet_1_1__leaf_net441),
    .S1(net968),
    .X(net705));
 sky130_fd_sc_hd__o2111ai_1 c732 (.A1(net685),
    .A2(net542),
    .B1(net937),
    .C1(net452),
    .D1(net319),
    .Y(net706));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net309),
    .A1(net512),
    .A2(net652),
    .A3(net633),
    .S0(net990),
    .S1(net885),
    .X(net707));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net687),
    .A1(net694),
    .A2(net999),
    .A3(net830),
    .S0(net849),
    .S1(net890),
    .X(net708));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(clknet_1_1__leaf_net679),
    .A1(clknet_1_1__leaf_net441),
    .A2(net309),
    .A3(net542),
    .S0(net698),
    .S1(net891),
    .X(net709));
 sky130_fd_sc_hd__mux4_4 c736 (.A0(net704),
    .A1(net672),
    .A2(clknet_1_1__leaf_net562),
    .A3(net150),
    .S0(net886),
    .S1(clknet_1_1__leaf_net892),
    .X(net710));
 sky130_fd_sc_hd__a2111oi_0 c737 (.A1(clknet_1_0__leaf_net665),
    .A2(net689),
    .B1(net684),
    .C1(net888),
    .D1(clknet_1_0__leaf_net892),
    .Y(net711));
 sky130_fd_sc_hd__mux4_2 c738 (.A0(net677),
    .A1(net708),
    .A2(net633),
    .A3(net652),
    .S0(clknet_1_1__leaf_net562),
    .S1(net886),
    .X(net712));
 sky130_fd_sc_hd__mux4_2 c739 (.A0(net706),
    .A1(clknet_1_0__leaf_net711),
    .A2(clknet_1_1__leaf_net665),
    .A3(clknet_1_0__leaf_net696),
    .S0(clknet_1_1__leaf_net562),
    .S1(net937),
    .X(net713));
 sky130_fd_sc_hd__nand2_4 c74 (.A(net42),
    .B(net938),
    .Y(net48));
 sky130_fd_sc_hd__mux4_2 c740 (.A0(net999),
    .A1(net710),
    .A2(net512),
    .A3(clknet_1_0__leaf_net711),
    .S0(net865),
    .S1(clknet_1_1__leaf_net892),
    .X(net714));
 sky130_fd_sc_hd__mux4_2 c741 (.A0(net672),
    .A1(net702),
    .A2(net988),
    .A3(net694),
    .S0(net886),
    .S1(clknet_1_0__leaf_net894),
    .X(net715));
 sky130_fd_sc_hd__mux4_4 c742 (.A0(net714),
    .A1(net695),
    .A2(clknet_1_0__leaf_net711),
    .A3(clknet_1_0__leaf_net715),
    .S0(clknet_1_0__leaf_net679),
    .S1(clknet_1_0__leaf_net894),
    .X(net716));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net452),
    .A1(net988),
    .A2(clknet_1_0__leaf_net711),
    .A3(net815),
    .S0(clknet_1_0__leaf_net892),
    .S1(net895),
    .X(net717));
 sky130_fd_sc_hd__mux4_2 c744 (.A0(net512),
    .A1(clknet_1_1__leaf_net715),
    .A2(net598),
    .A3(clknet_1_1__leaf_net711),
    .S0(clknet_1_0__leaf_net894),
    .S1(net895),
    .X(net718));
 sky130_fd_sc_hd__mux4_4 c745 (.A0(net703),
    .A1(clknet_1_0__leaf_net715),
    .A2(clknet_1_0__leaf_net711),
    .A3(net865),
    .S0(clknet_1_1__leaf_net892),
    .S1(clknet_1_0__leaf_net894),
    .X(net719));
 sky130_fd_sc_hd__mux4_2 c746 (.A0(net719),
    .A1(net717),
    .A2(clknet_1_0__leaf_net711),
    .A3(net599),
    .S0(net685),
    .S1(clknet_1_1__leaf_net894),
    .X(net720));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net319),
    .A1(net718),
    .A2(net542),
    .A3(clknet_1_1__leaf_net715),
    .S0(net893),
    .S1(net898),
    .X(net721));
 sky130_fd_sc_hd__mux4_4 c748 (.A0(clknet_1_1__leaf_net711),
    .A1(net985),
    .A2(clknet_1_1__leaf_net696),
    .A3(net1037),
    .S0(net849),
    .S1(net897),
    .X(net722));
 sky130_fd_sc_hd__mux4_4 c749 (.A0(net619),
    .A1(net56),
    .A2(net998),
    .A3(net869),
    .S0(net896),
    .S1(net897),
    .X(net723));
 sky130_fd_sc_hd__or2b_1 c75 (.A(net35),
    .B_N(net48),
    .X(net49));
 sky130_fd_sc_hd__mux4_2 c750 (.A0(clknet_1_1__leaf_net346),
    .A1(net937),
    .A2(net796),
    .A3(net867),
    .S0(clknet_1_1__leaf_net894),
    .S1(net896),
    .X(net724));
 sky130_fd_sc_hd__mux4_4 c751 (.A0(clknet_1_0__leaf_net724),
    .A1(net869),
    .A2(net890),
    .A3(net898),
    .S0(net900),
    .S1(net901),
    .X(net725));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(clknet_1_0__leaf_net724),
    .A1(net725),
    .A2(clknet_1_1__leaf_net711),
    .A3(net204),
    .S0(net869),
    .S1(net890),
    .X(net726));
 sky130_fd_sc_hd__mux4_4 c753 (.A0(net988),
    .A1(clknet_1_1__leaf_net674),
    .A2(clknet_1_0__leaf_net696),
    .A3(net890),
    .S0(clknet_1_1__leaf_net894),
    .S1(net896),
    .X(net727));
 sky130_fd_sc_hd__mux4_2 c754 (.A0(net617),
    .A1(net204),
    .A2(net968),
    .A3(clknet_1_1__leaf_net346),
    .S0(net179),
    .S1(clknet_1_1__leaf_net464),
    .X(net728));
 sky130_fd_sc_hd__mux4_4 c755 (.A0(net208),
    .A1(net998),
    .A2(clknet_1_1__leaf_net674),
    .A3(clknet_1_1__leaf_net894),
    .S0(net898),
    .S1(net901),
    .X(net729));
 sky130_fd_sc_hd__mux4_4 c756 (.A0(net625),
    .A1(clknet_1_1__leaf_net665),
    .A2(net726),
    .A3(net699),
    .S0(net179),
    .S1(net869),
    .X(net730));
 sky130_fd_sc_hd__mux4_4 c757 (.A0(net985),
    .A1(clknet_1_1__leaf_net464),
    .A2(clknet_1_1__leaf_net674),
    .A3(net901),
    .S0(net902),
    .S1(net903),
    .X(net731));
 sky130_fd_sc_hd__mux4_2 c758 (.A0(net563),
    .A1(clknet_1_1__leaf_net696),
    .A2(net937),
    .A3(clknet_1_1__leaf_net728),
    .S0(net902),
    .S1(net903),
    .X(net732));
 sky130_fd_sc_hd__mux4_2 c759 (.A0(clknet_1_1__leaf_net486),
    .A1(net699),
    .A2(net886),
    .A3(net890),
    .S0(net899),
    .S1(net902),
    .X(net733));
 sky130_fd_sc_hd__and2b_2 c76 (.A_N(net19),
    .B(net29),
    .X(net50));
 sky130_fd_sc_hd__sdfbbp_1 c760 (.CLK(clknet_4_13_0_clk),
    .D(net652),
    .RESET_B(clknet_1_1__leaf_net724),
    .SCD(clknet_1_0__leaf_net728),
    .SCE(net56),
    .SET_B(net806),
    .Q(net734));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(clknet_1_1__leaf_net665),
    .A1(clknet_1_1__leaf_net724),
    .A2(net903),
    .A3(net904),
    .S0(net905),
    .S1(net906),
    .X(net735));
 sky130_fd_sc_hd__mux4_2 c762 (.A0(net690),
    .A1(clknet_1_0__leaf_net728),
    .A2(net734),
    .A3(net735),
    .S0(clknet_1_1__leaf_net346),
    .S1(net208));
 sky130_fd_sc_hd__or3b_1 c77 (.A(net26),
    .B(net42),
    .C_N(net48),
    .X(net51));
 sky130_fd_sc_hd__nand2b_2 c78 (.A_N(net0),
    .B(net47),
    .Y(net52));
 sky130_fd_sc_hd__nand2b_1 c79 (.A_N(net50),
    .B(net51),
    .Y(net53));
 sky130_fd_sc_hd__buf_6 c80 (.A(net794),
    .X(net54));
 sky130_fd_sc_hd__nor2_4 c81 (.A(net50),
    .B(net45),
    .Y(net55));
 sky130_fd_sc_hd__buf_4 c82 (.A(net794),
    .X(net56));
 sky130_fd_sc_hd__nor3b_1 c83 (.A(net47),
    .B(net51),
    .C_N(net999),
    .Y(net57));
 sky130_fd_sc_hd__nor3b_1 c84 (.A(net21),
    .B(net50),
    .C_N(net49),
    .Y(net58));
 sky130_fd_sc_hd__sdfbbn_1 c85 (.CLK_N(clknet_4_8_0_clk),
    .D(net49),
    .RESET_B(net58),
    .SCD(net47),
    .SCE(net999),
    .SET_B(net48),
    .Q(net60),
    .Q_N(net59));
 sky130_fd_sc_hd__clkbuf_2 c86 (.A(net828),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 c87 (.A(net916),
    .X(net62));
 sky130_fd_sc_hd__and2b_1 c88 (.A_N(net33),
    .B(net1004),
    .X(net63));
 sky130_fd_sc_hd__or2_1 c89 (.A(net999),
    .B(net29),
    .X(net64));
 sky130_fd_sc_hd__or3b_2 c90 (.A(net51),
    .B(net1004),
    .C_N(net982),
    .X(net65));
 sky130_fd_sc_hd__nand2_1 c91 (.A(net64),
    .B(net60),
    .Y(net66));
 sky130_fd_sc_hd__buf_1 c92 (.A(net918),
    .X(net67));
 sky130_fd_sc_hd__nor3b_1 c93 (.A(net935),
    .B(net64),
    .C_N(net18),
    .Y(net68));
 sky130_fd_sc_hd__and2_1 c94 (.A(net63),
    .B(net64),
    .X(net69));
 sky130_fd_sc_hd__or4bb_1 c95 (.A(net986),
    .B(net29),
    .C_N(net935),
    .D_N(net48),
    .X(net70));
 sky130_fd_sc_hd__nor2b_2 c96 (.A(net45),
    .B_N(net59),
    .Y(net71));
 sky130_fd_sc_hd__nor2_1 c97 (.A(net71),
    .B(net986),
    .Y(net72));
 sky130_fd_sc_hd__nand2b_2 c98 (.A_N(net27),
    .B(net63),
    .Y(net73));
 sky130_fd_sc_hd__nor2_1 c99 (.A(net60),
    .B(net66),
    .Y(net74));
 sky130_fd_sc_hd__sdfbbn_1 merge763 (.CLK_N(clknet_4_9_0_clk),
    .D(net337),
    .RESET_B(net195),
    .SCD(net340),
    .SCE(net158),
    .SET_B(clknet_1_0__leaf_net210),
    .Q(net737),
    .Q_N(net736));
 sky130_fd_sc_hd__buf_16 merge764 (.A(net794),
    .X(net738));
 sky130_fd_sc_hd__sdfbbn_1 merge765 (.CLK_N(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net641),
    .RESET_B(net389),
    .SCD(net654),
    .SCE(net555),
    .SET_B(net1042),
    .Q(net740),
    .Q_N(net739));
 sky130_fd_sc_hd__sdfrtp_4 merge766 (.CLK(clknet_4_8_0_clk),
    .D(net1034),
    .RESET_B(net65),
    .SCD(net983),
    .SCE(net195),
    .Q(net741));
 sky130_fd_sc_hd__inv_4 merge767 (.A(net920),
    .Y(net742));
 sky130_fd_sc_hd__sdfbbp_1 merge768 (.CLK(clknet_4_6_0_clk),
    .D(net325),
    .RESET_B(net423),
    .SCD(clknet_1_1__leaf_net583),
    .SCE(net142),
    .SET_B(net405),
    .Q(net744),
    .Q_N(net743));
 sky130_fd_sc_hd__or4bb_1 merge769 (.A(net76),
    .B(net45),
    .C_N(net69),
    .D_N(net74),
    .X(net745));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(net14),
    .A1(net158),
    .A2(net927),
    .A3(net34),
    .S0(net159),
    .S1(net163),
    .X(net746));
 sky130_fd_sc_hd__a2111oi_1 merge771 (.A1(net399),
    .A2(net407),
    .B1(net270),
    .C1(net133),
    .D1(net278),
    .Y(net747));
 sky130_fd_sc_hd__or4bb_2 merge772 (.A(net278),
    .B(net260),
    .C_N(clknet_1_1__leaf_net532),
    .D_N(net422),
    .X(net748));
 sky130_fd_sc_hd__or4bb_1 merge773 (.A(net265),
    .B(net381),
    .C_N(net382),
    .D_N(net112),
    .X(net749));
 sky130_fd_sc_hd__mux4_2 merge774 (.A0(net17),
    .A1(net386),
    .A2(net428),
    .A3(net1000),
    .S0(clknet_1_0__leaf_net430),
    .S1(net1003),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd1_1 merge775 (.A(net917),
    .X(net751));
 sky130_fd_sc_hd__mux4_4 merge776 (.A0(net630),
    .A1(net513),
    .A2(clknet_1_1__leaf_net534),
    .A3(clknet_1_1__leaf_net639),
    .S0(net642),
    .S1(net643),
    .X(net752));
 sky130_fd_sc_hd__sdfrtp_1 merge777 (.CLK(clknet_4_2_0_clk),
    .D(net12),
    .RESET_B(net163),
    .SCE(net288),
    .Q(net289));
 sky130_fd_sc_hd__sdfsbp_1 merge778 (.CLK(clknet_4_10_0_clk),
    .D(net193),
    .SCD(net974),
    .SCE(net100),
    .SET_B(net979),
    .Q(net755),
    .Q_N(net754));
 sky130_fd_sc_hd__sdfbbn_1 merge779 (.CLK_N(clknet_4_10_0_clk),
    .D(net84),
    .RESET_B(net979),
    .SCD(clknet_1_0__leaf_net83),
    .SCE(net974),
    .SET_B(net983),
    .Q(net757),
    .Q_N(net756));
 sky130_fd_sc_hd__sdfsbp_1 merge780 (.CLK(clknet_4_9_0_clk),
    .D(net195),
    .SCD(net980),
    .SCE(net181),
    .SET_B(net323),
    .Q(net759),
    .Q_N(net758));
 sky130_fd_sc_hd__inv_2 merge781 (.A(net829),
    .Y(net760));
 sky130_fd_sc_hd__or4bb_1 merge782 (.A(net451),
    .B(net316),
    .C_N(net296),
    .D_N(net298),
    .X(net761));
 sky130_fd_sc_hd__or4bb_1 merge783 (.A(net31),
    .B(net180),
    .C_N(net293),
    .D_N(net978),
    .X(net762));
 sky130_fd_sc_hd__or4bb_2 merge784 (.A(net53),
    .B(net27),
    .C_N(net979),
    .D_N(clknet_1_0__leaf_net201),
    .X(net763));
 sky130_fd_sc_hd__mux4_4 merge785 (.A0(net550),
    .A1(net538),
    .A2(net542),
    .A3(net422),
    .S0(net544),
    .S1(net547),
    .X(net764));
 sky130_fd_sc_hd__sdfstp_1 merge786 (.CLK(clknet_4_3_0_clk),
    .D(net255),
    .SCD(net288),
    .SCE(net327),
    .SET_B(net934),
    .Q(net765));
 sky130_fd_sc_hd__mux4_2 merge787 (.A0(clknet_1_1__leaf_net664),
    .A1(net676),
    .A2(net549),
    .A3(net386),
    .S0(net558),
    .S1(net889),
    .X(net766));
 sky130_fd_sc_hd__mux4_2 merge788 (.A0(net301),
    .A1(net291),
    .A2(net988),
    .A3(clknet_1_0__leaf_net81),
    .S0(clknet_1_0__leaf_net339),
    .S1(net1002),
    .X(net767));
 sky130_fd_sc_hd__sdfstp_1 merge789 (.CLK(clknet_4_11_0_clk),
    .D(net228),
    .SCD(net1028),
    .SCE(net974),
    .SET_B(clknet_1_1__leaf_net227),
    .Q(net768));
 sky130_fd_sc_hd__sdfstp_1 merge790 (.CLK(clknet_4_0_0_clk),
    .D(net383),
    .SCD(net516),
    .SCE(net393),
    .SET_B(net382),
    .Q(net769));
 sky130_fd_sc_hd__a2111oi_1 merge791 (.A1(net42),
    .A2(net53),
    .B1(net180),
    .C1(net154),
    .D1(net188),
    .Y(net770));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net163),
    .A1(net166),
    .A2(net253),
    .A3(net272),
    .S0(net280),
    .S1(net811),
    .X(net771));
 sky130_fd_sc_hd__mux4_2 merge793 (.A0(clknet_1_0__leaf_net657),
    .A1(net653),
    .A2(clknet_1_1__leaf_net641),
    .A3(net154),
    .S0(net407),
    .S1(net251),
    .X(net772));
 sky130_fd_sc_hd__mux4_4 merge794 (.A0(net65),
    .A1(net153),
    .A2(net79),
    .A3(net73),
    .S0(clknet_1_0__leaf_net227),
    .S1(clknet_1_0__leaf_net214),
    .X(net773));
 sky130_fd_sc_hd__buf_1 merge795 (.A(net919),
    .X(net774));
 sky130_fd_sc_hd__o2111ai_1 merge796 (.A1(net157),
    .A2(net184),
    .B1(net195),
    .C1(net46),
    .D1(net970),
    .Y(net775));
 sky130_fd_sc_hd__buf_6 merge797 (.A(net829),
    .X(net776));
 sky130_fd_sc_hd__mux4_1 merge798 (.A0(net996),
    .A1(net406),
    .A2(net519),
    .A3(net643),
    .S0(net403),
    .S1(net846),
    .X(net777));
 sky130_fd_sc_hd__mux4_1 merge799 (.A0(net170),
    .A1(net168),
    .A2(net174),
    .A3(net58),
    .S0(net53),
    .S1(net50),
    .X(net778));
 sky130_fd_sc_hd__mux4_1 merge800 (.A0(net383),
    .A1(net123),
    .A2(net942),
    .A3(net385),
    .S0(net382),
    .S1(net391),
    .X(net779));
 sky130_fd_sc_hd__mux4_2 merge801 (.A0(net398),
    .A1(net382),
    .A2(net385),
    .A3(net443),
    .S0(clknet_1_0__leaf_net822),
    .S1(clknet_1_0__leaf_net967),
    .X(net780));
 sky130_fd_sc_hd__mux4_4 merge802 (.A0(net58),
    .A1(net59),
    .A2(net61),
    .A3(net213),
    .S0(net73),
    .S1(net1002),
    .X(net781));
 sky130_fd_sc_hd__mux4_4 merge803 (.A0(net62),
    .A1(net65),
    .A2(net934),
    .A3(net41),
    .S0(net44),
    .S1(net933),
    .X(net782));
 sky130_fd_sc_hd__mux4_1 merge804 (.A0(net942),
    .A1(net386),
    .A2(net264),
    .A3(net932),
    .S0(net517),
    .S1(net515),
    .X(net783));
 sky130_fd_sc_hd__sdfbbn_1 merge805 (.CLK_N(clknet_4_3_0_clk),
    .D(net282),
    .RESET_B(net386),
    .SCD(net260),
    .SCE(net428),
    .SET_B(clknet_1_0__leaf_net972),
    .Q(net785),
    .Q_N(net784));
 sky130_fd_sc_hd__sdfbbp_1 merge806 (.CLK(clknet_4_0_0_clk),
    .D(net407),
    .RESET_B(net151),
    .SCD(net410),
    .SCE(net996),
    .SET_B(net417),
    .Q(net787),
    .Q_N(net786));
 sky130_fd_sc_hd__mux4_1 merge807 (.A0(net1),
    .A1(net405),
    .A2(net407),
    .A3(net280),
    .S0(net403),
    .S1(net414),
    .X(net788));
 sky130_fd_sc_hd__mux4_1 merge808 (.A0(net406),
    .A1(net415),
    .A2(net252),
    .A3(net543),
    .S0(net546),
    .S1(net975),
    .X(net789));
 sky130_fd_sc_hd__dfrbp_1 merge809 (.CLK(clknet_4_10_0_clk),
    .D(net102),
    .RESET_B(net109),
    .Q(net791),
    .Q_N(net790));
 sky130_fd_sc_hd__dfrbp_1 merge810 (.CLK(clknet_4_9_0_clk),
    .D(net326),
    .RESET_B(net333),
    .Q(net793),
    .Q_N(net792));
 sky130_fd_sc_hd__dfrtn_1 merge811 (.CLK_N(clknet_4_8_0_clk),
    .D(net763),
    .RESET_B(net1060),
    .Q(net794));
 sky130_fd_sc_hd__dfrtp_1 merge812 (.CLK(clknet_4_9_0_clk),
    .D(net211),
    .RESET_B(net217),
    .Q(net795));
 sky130_fd_sc_hd__dfrtp_1 merge813 (.CLK(clknet_4_12_0_clk),
    .D(net470),
    .RESET_B(net477),
    .Q(net796));
 sky130_fd_sc_hd__dfrtp_2 merge814 (.CLK(clknet_4_11_0_clk),
    .D(net235),
    .RESET_B(net242),
    .Q(net797));
 sky130_fd_sc_hd__dfsbp_1 merge815 (.CLK(clknet_4_11_0_clk),
    .D(net357),
    .SET_B(net362),
    .Q(net799),
    .Q_N(net798));
 sky130_fd_sc_hd__dfsbp_1 merge816 (.CLK(clknet_4_5_0_clk),
    .D(net648),
    .SET_B(net667),
    .Q(net801),
    .Q_N(net800));
 sky130_fd_sc_hd__dfstp_1 merge817 (.CLK(clknet_4_6_0_clk),
    .D(net586),
    .SET_B(net597),
    .Q(net802));
 sky130_fd_sc_hd__dfstp_2 merge818 (.CLK(clknet_4_9_0_clk),
    .D(net762),
    .SET_B(net775),
    .Q(net803));
 sky130_fd_sc_hd__and2b_1 merge819 (.A_N(net680),
    .B(net683),
    .X(net804));
 sky130_fd_sc_hd__dfstp_1 merge820 (.CLK(clknet_4_1_0_clk),
    .D(net530),
    .SET_B(net535),
    .Q(net805));
 sky130_fd_sc_hd__dlrbn_1 merge821 (.D(net722),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net730),
    .Q(net806));
 sky130_fd_sc_hd__dlrbn_1 merge822 (.D(net495),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net496),
    .Q(net807),
    .Q_N(net958));
 sky130_fd_sc_hd__dlrbp_1 merge823 (.D(net177),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net746),
    .Q(net809),
    .Q_N(net808));
 sky130_fd_sc_hd__dlrbp_1 merge824 (.D(net275),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net276),
    .Q(net811),
    .Q_N(net810));
 sky130_fd_sc_hd__dlrtn_1 merge825 (.D(net603),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net605),
    .Q(net812));
 sky130_fd_sc_hd__dlrtn_1 merge826 (.D(net424),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net973),
    .Q(net813));
 sky130_fd_sc_hd__dlrtn_1 merge827 (.D(net303),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net310),
    .Q(net814));
 sky130_fd_sc_hd__dlrtp_1 merge828 (.D(net700),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net701),
    .Q(net815));
 sky130_fd_sc_hd__dlrtp_1 merge829 (.D(net453),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net761),
    .Q(net816));
 sky130_fd_sc_hd__dlrtp_1 merge830 (.D(net748),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net764),
    .Q(net817));
 sky130_fd_sc_hd__edfxbp_1 merge831 (.CLK(clknet_4_9_0_clk),
    .D(net342),
    .DE(net347),
    .Q(net819),
    .Q_N(net818));
 sky130_fd_sc_hd__edfxtp_1 merge832 (.CLK(clknet_4_5_0_clk),
    .D(net646),
    .DE(net752),
    .Q(net820));
 sky130_fd_sc_hd__sdlclkp_1 merge833 (.CLK(clknet_4_6_0_clk),
    .GATE(net559),
    .SCE(net565),
    .GCLK(net821));
 sky130_fd_sc_hd__sdlclkp_2 merge834 (.CLK(clknet_4_3_0_clk),
    .GATE(net436),
    .SCE(net446),
    .GCLK(net822));
 sky130_fd_sc_hd__sdlclkp_4 merge835 (.CLK(clknet_4_8_0_clk),
    .GATE(net80),
    .SCE(net745),
    .GCLK(net823));
 sky130_fd_sc_hd__dfrbp_2 merge836 (.CLK(clknet_4_0_0_clk),
    .D(net402),
    .RESET_B(net749),
    .Q(net825),
    .Q_N(net824));
 sky130_fd_sc_hd__dfrbp_1 merge837 (.CLK(clknet_4_15_0_clk),
    .D(net479),
    .RESET_B(net511),
    .Q(net827),
    .Q_N(net826));
 sky130_fd_sc_hd__dfrtn_1 merge838 (.CLK_N(clknet_4_8_0_clk),
    .D(net220),
    .RESET_B(net778),
    .Q(net828));
 sky130_fd_sc_hd__dfrtp_4 merge839 (.CLK(clknet_4_0_0_clk),
    .D(net779),
    .RESET_B(net780),
    .Q(net829));
 sky130_fd_sc_hd__dfrtp_1 merge840 (.CLK(clknet_4_15_0_clk),
    .D(net480),
    .RESET_B(net509),
    .Q(net963));
 sky130_fd_sc_hd__dfrtp_1 merge841 (.CLK(clknet_4_5_0_clk),
    .D(net697),
    .RESET_B(net804),
    .Q(net830));
 sky130_fd_sc_hd__dfsbp_1 merge842 (.CLK(clknet_4_14_0_clk),
    .D(net481),
    .SET_B(net508),
    .Q(net831),
    .Q_N(net948));
 sky130_fd_sc_hd__dfxbp_1 s843 (.CLK(clknet_4_8_0_clk),
    .D(net82),
    .Q(net833),
    .Q_N(net832));
 sky130_fd_sc_hd__dfxbp_1 s844 (.CLK(clknet_4_11_0_clk),
    .D(net108),
    .Q(net835),
    .Q_N(net834));
 sky130_fd_sc_hd__dfxtp_2 s845 (.CLK(clknet_4_11_0_clk),
    .D(net110),
    .Q(net836));
 sky130_fd_sc_hd__dfxtp_1 s846 (.CLK(clknet_4_2_0_clk),
    .D(net171),
    .Q(net837));
 sky130_fd_sc_hd__dfxtp_1 s847 (.CLK(clknet_4_2_0_clk),
    .D(net176),
    .Q(net838));
 sky130_fd_sc_hd__dlclkp_1 s848 (.CLK(clknet_4_8_0_clk),
    .GATE(net219),
    .GCLK(net839));
 sky130_fd_sc_hd__dlclkp_2 s849 (.CLK(clknet_4_10_0_clk),
    .GATE(net236),
    .GCLK(net840));
 sky130_fd_sc_hd__dlclkp_4 s850 (.CLK(clknet_4_14_0_clk),
    .GATE(net243),
    .GCLK(net841));
 sky130_fd_sc_hd__dlxbn_1 s851 (.D(net244),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net843),
    .Q_N(net842));
 sky130_fd_sc_hd__dlxbn_2 s852 (.D(net285),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net845),
    .Q_N(net844));
 sky130_fd_sc_hd__dlxbp_1 s853 (.D(net286),
    .GATE(clknet_4_1_0_clk),
    .Q(net847),
    .Q_N(net846));
 sky130_fd_sc_hd__dlxtn_2 s854 (.D(net305),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net971));
 sky130_fd_sc_hd__dlxtn_1 s855 (.D(net334),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net848));
 sky130_fd_sc_hd__dlxtn_2 s856 (.D(net335),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net849));
 sky130_fd_sc_hd__dlxtp_1 s857 (.D(net353),
    .GATE(clknet_4_9_0_clk),
    .Q(net850));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s858 (.D(net368),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net851));
 sky130_fd_sc_hd__dfxbp_1 s859 (.CLK(clknet_4_11_0_clk),
    .D(net369),
    .Q(net853),
    .Q_N(net852));
 sky130_fd_sc_hd__dfxbp_1 s860 (.CLK(clknet_4_11_0_clk),
    .D(net371),
    .Q(net854));
 sky130_fd_sc_hd__dfxtp_1 s861 (.CLK(clknet_4_11_0_clk),
    .D(net374),
    .Q(net855));
 sky130_fd_sc_hd__dfxtp_1 s862 (.CLK(clknet_4_14_0_clk),
    .D(net375),
    .Q(net856));
 sky130_fd_sc_hd__dfxtp_1 s863 (.CLK(clknet_4_14_0_clk),
    .D(net378),
    .Q(net857));
 sky130_fd_sc_hd__dlclkp_1 s864 (.CLK(clknet_4_14_0_clk),
    .GATE(net380),
    .GCLK(net858));
 sky130_fd_sc_hd__dlclkp_2 s865 (.CLK(clknet_4_3_0_clk),
    .GATE(net437),
    .GCLK(net972));
 sky130_fd_sc_hd__dlclkp_4 s866 (.CLK(clknet_4_3_0_clk),
    .GATE(net438),
    .GCLK(net967));
 sky130_fd_sc_hd__dlxbn_1 s867 (.D(net445),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net860),
    .Q_N(net859));
 sky130_fd_sc_hd__dlxbn_1 s868 (.D(net447),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net862),
    .Q_N(net861));
 sky130_fd_sc_hd__dlxbp_1 s869 (.D(net462),
    .GATE(clknet_4_12_0_clk),
    .Q(net864),
    .Q_N(net863));
 sky130_fd_sc_hd__dlxtn_1 s870 (.D(net465),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net865));
 sky130_fd_sc_hd__dlxtn_1 s871 (.D(net468),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net866));
 sky130_fd_sc_hd__dlxtn_2 s872 (.D(net469),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net867));
 sky130_fd_sc_hd__dlxtp_1 s873 (.D(net482),
    .GATE(clknet_4_12_0_clk),
    .Q(net868));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s874 (.D(net494),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net869));
 sky130_fd_sc_hd__dfxbp_1 s875 (.CLK(clknet_4_15_0_clk),
    .D(net497),
    .Q(net870));
 sky130_fd_sc_hd__dfxbp_1 s876 (.CLK(clknet_4_14_0_clk),
    .D(net500),
    .Q(net872),
    .Q_N(net871));
 sky130_fd_sc_hd__dfxtp_1 s877 (.CLK(clknet_4_15_0_clk),
    .D(net503),
    .Q(net962));
 sky130_fd_sc_hd__dfxtp_2 s878 (.CLK(clknet_4_15_0_clk),
    .D(net505),
    .Q(net873));
 sky130_fd_sc_hd__dfxtp_1 s879 (.CLK(clknet_4_15_0_clk),
    .D(net506),
    .Q(net874));
 sky130_fd_sc_hd__dlclkp_1 s880 (.CLK(clknet_4_15_0_clk),
    .GATE(net507),
    .GCLK(net964));
 sky130_fd_sc_hd__dlclkp_2 s881 (.CLK(clknet_4_15_0_clk),
    .GATE(net510),
    .GCLK(net875));
 sky130_fd_sc_hd__dlclkp_4 s882 (.CLK(clknet_4_1_0_clk),
    .GATE(net531),
    .GCLK(net876));
 sky130_fd_sc_hd__dlxbn_1 s883 (.D(net569),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net878),
    .Q_N(net877));
 sky130_fd_sc_hd__dlxbn_1 s884 (.D(net575),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net880),
    .Q_N(net879));
 sky130_fd_sc_hd__dlxbp_1 s885 (.D(net594),
    .GATE(clknet_4_7_0_clk),
    .Q(net882),
    .Q_N(net881));
 sky130_fd_sc_hd__dlxtn_1 s886 (.D(net595),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net883));
 sky130_fd_sc_hd__dlxtn_2 s887 (.D(net596),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net952));
 sky130_fd_sc_hd__dlxtn_1 s888 (.D(net600),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net955));
 sky130_fd_sc_hd__dlxtp_1 s889 (.D(net604),
    .GATE(clknet_4_13_0_clk),
    .Q(net961));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s890 (.D(net622),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net884));
 sky130_fd_sc_hd__dfxbp_2 s891 (.CLK(clknet_4_5_0_clk),
    .D(net647),
    .Q(net886),
    .Q_N(net885));
 sky130_fd_sc_hd__dfxbp_1 s892 (.CLK(clknet_4_5_0_clk),
    .D(net670),
    .Q(net888),
    .Q_N(net887));
 sky130_fd_sc_hd__dfxtp_2 s893 (.CLK(clknet_4_5_0_clk),
    .D(net686),
    .Q(net889));
 sky130_fd_sc_hd__dfxtp_1 s894 (.CLK(clknet_4_7_0_clk),
    .D(net705),
    .Q(net890));
 sky130_fd_sc_hd__dfxtp_1 s895 (.CLK(clknet_4_5_0_clk),
    .D(net707),
    .Q(net891));
 sky130_fd_sc_hd__dlclkp_1 s896 (.CLK(clknet_4_7_0_clk),
    .GATE(net709),
    .GCLK(net892));
 sky130_fd_sc_hd__dlclkp_2 s897 (.CLK(clknet_4_7_0_clk),
    .GATE(net712),
    .GCLK(net893));
 sky130_fd_sc_hd__dlclkp_4 s898 (.CLK(clknet_4_7_0_clk),
    .GATE(net713),
    .GCLK(net894));
 sky130_fd_sc_hd__dlxbn_1 s899 (.D(net716),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net896),
    .Q_N(net895));
 sky130_fd_sc_hd__dlxbn_1 s900 (.D(net720),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net898),
    .Q_N(net897));
 sky130_fd_sc_hd__dlxbp_1 s901 (.D(net721),
    .GATE(clknet_4_7_0_clk),
    .Q(net900),
    .Q_N(net899));
 sky130_fd_sc_hd__dlxtn_1 s902 (.D(net723),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net901));
 sky130_fd_sc_hd__dlxtn_1 s903 (.D(net727),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net902));
 sky130_fd_sc_hd__dlxtn_1 s904 (.D(net729),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net903));
 sky130_fd_sc_hd__dlxtp_1 s905 (.D(net731),
    .GATE(clknet_4_13_0_clk),
    .Q(net904));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s906 (.D(net732),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net905));
 sky130_fd_sc_hd__dfxbp_1 s907 (.CLK(clknet_4_13_0_clk),
    .D(net733),
    .Q(net906));
 sky130_fd_sc_hd__dfxbp_1 s908 (.CLK(clknet_4_6_0_clk),
    .D(net750),
    .Q(net908),
    .Q_N(net907));
 sky130_fd_sc_hd__dfxtp_1 s909 (.CLK(clknet_4_4_0_clk),
    .D(net766),
    .Q(net909));
 sky130_fd_sc_hd__dfxtp_1 s910 (.CLK(clknet_4_9_0_clk),
    .D(net767),
    .Q(net910));
 sky130_fd_sc_hd__dfxtp_1 s911 (.CLK(clknet_4_2_0_clk),
    .D(net771),
    .Q(net911));
 sky130_fd_sc_hd__dlclkp_1 s912 (.CLK(clknet_4_1_0_clk),
    .GATE(net772),
    .GCLK(net912));
 sky130_fd_sc_hd__dlclkp_2 s913 (.CLK(clknet_4_11_0_clk),
    .GATE(net773),
    .GCLK(net913));
 sky130_fd_sc_hd__dlclkp_4 s914 (.CLK(clknet_4_0_0_clk),
    .GATE(net777),
    .GCLK(net914));
 sky130_fd_sc_hd__dlxbn_1 s915 (.D(net781),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net916),
    .Q_N(net915));
 sky130_fd_sc_hd__dlxbn_1 s916 (.D(net782),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net918),
    .Q_N(net917));
 sky130_fd_sc_hd__dlxbp_1 s917 (.D(net783),
    .GATE(clknet_4_1_0_clk),
    .Q(net920),
    .Q_N(net919));
 sky130_fd_sc_hd__dlxtn_1 s918 (.D(net788),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net921));
 sky130_fd_sc_hd__dlxtn_1 s919 (.D(net789),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net922));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_8 input2 (.A(in1),
    .X(net924));
 sky130_fd_sc_hd__buf_2 input3 (.A(in10),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(in11),
    .X(net926));
 sky130_fd_sc_hd__buf_2 input5 (.A(in12),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_8 input6 (.A(in13),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in14),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in15),
    .X(net930));
 sky130_fd_sc_hd__buf_2 input9 (.A(in16),
    .X(net931));
 sky130_fd_sc_hd__buf_1 input10 (.A(in17),
    .X(net932));
 sky130_fd_sc_hd__buf_1 input11 (.A(in18),
    .X(net933));
 sky130_fd_sc_hd__buf_4 input12 (.A(in19),
    .X(net934));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(in2),
    .X(net935));
 sky130_fd_sc_hd__buf_2 input14 (.A(in20),
    .X(net936));
 sky130_fd_sc_hd__buf_12 input15 (.A(in21),
    .X(net937));
 sky130_fd_sc_hd__buf_2 input16 (.A(in22),
    .X(net938));
 sky130_fd_sc_hd__buf_2 input17 (.A(in23),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in24),
    .X(net940));
 sky130_fd_sc_hd__buf_2 input19 (.A(in3),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in4),
    .X(net942));
 sky130_fd_sc_hd__buf_6 input21 (.A(in5),
    .X(net943));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(in6),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in7),
    .X(net945));
 sky130_fd_sc_hd__buf_1 input24 (.A(in8),
    .X(net946));
 sky130_fd_sc_hd__buf_4 input25 (.A(in9),
    .X(net947));
 sky130_fd_sc_hd__buf_2 output26 (.A(net948),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output27 (.A(net949),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output28 (.A(net950),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output29 (.A(net951),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net952),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output31 (.A(net953),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output32 (.A(net954),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output33 (.A(net955),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net956),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(clknet_1_1__leaf_net957),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output36 (.A(net958),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output37 (.A(net981),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output38 (.A(net960),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output39 (.A(net961),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output40 (.A(net962),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output41 (.A(net963),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net964),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net965),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output44 (.A(net966),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(clknet_1_1__leaf_net967),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output46 (.A(net968),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output47 (.A(net969),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net1009),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output49 (.A(net971),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(clknet_1_1__leaf_net972),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_1 wire51 (.A(net747),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_2 wire52 (.A(net57),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(net423),
    .X(net975));
 sky130_fd_sc_hd__buf_1 max_cap54 (.A(net336),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_1 max_cap55 (.A(net317),
    .X(net977));
 sky130_fd_sc_hd__buf_1 max_cap56 (.A(net165),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net79),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(net959),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net38),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout61 (.A(net38),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_2 max_cap62 (.A(net290),
    .X(net984));
 sky130_fd_sc_hd__buf_4 fanout63 (.A(net150),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_2 max_cap64 (.A(net68),
    .X(net986));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(net208),
    .X(net987));
 sky130_fd_sc_hd__buf_4 fanout66 (.A(net179),
    .X(net988));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap67 (.A(net991),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_2 max_cap68 (.A(net991),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_2 wire69 (.A(net992),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_2 max_cap70 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_2 max_cap71 (.A(net16),
    .X(net993));
 sky130_fd_sc_hd__clkbuf_2 wire72 (.A(net995),
    .X(net994));
 sky130_fd_sc_hd__buf_6 wire73 (.A(net128),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_2 max_cap74 (.A(net127),
    .X(net996));
 sky130_fd_sc_hd__buf_6 fanout75 (.A(net9),
    .X(net997));
 sky130_fd_sc_hd__buf_4 max_cap76 (.A(net5),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_4 fanout77 (.A(net56),
    .X(net999));
 sky130_fd_sc_hd__buf_4 fanout78 (.A(net953),
    .X(net1000));
 sky130_fd_sc_hd__buf_4 fanout79 (.A(net971),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(net838),
    .X(net1002));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(net838),
    .X(net1003));
 sky130_fd_sc_hd__buf_2 fanout82 (.A(net39),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(net951),
    .X(net1005));
 sky130_fd_sc_hd__buf_8 fanout84 (.A(net1007),
    .X(net1006));
 sky130_fd_sc_hd__buf_12 fanout85 (.A(net1008),
    .X(net1007));
 sky130_fd_sc_hd__buf_12 fanout86 (.A(net113),
    .X(net1008));
 sky130_fd_sc_hd__inv_16 c104_1 (.A(clknet_1_0__leaf_net823),
    .Y(net1009));
 sky130_fd_sc_hd__inv_16 net999_2 (.A(clknet_1_1__leaf_net823),
    .Y(net1010));
 sky130_fd_sc_hd__inv_16 net999_3 (.A(clknet_1_1__leaf_net823),
    .Y(net1011));
 sky130_fd_sc_hd__inv_16 net999_4 (.A(clknet_1_1__leaf_net823),
    .Y(net1012));
 sky130_fd_sc_hd__inv_16 net999_5 (.A(clknet_1_1__leaf_net823),
    .Y(net1013));
 sky130_fd_sc_hd__inv_16 net999_6 (.A(clknet_1_1__leaf_net823),
    .Y(net1014));
 sky130_fd_sc_hd__inv_16 net999_7 (.A(clknet_1_0__leaf_net823),
    .Y(net1015));
 sky130_fd_sc_hd__inv_16 net999_8 (.A(clknet_1_0__leaf_net823),
    .Y(net1016));
 sky130_fd_sc_hd__inv_16 net999_9 (.A(clknet_1_0__leaf_net823),
    .Y(net1017));
 sky130_fd_sc_hd__inv_16 net999_10 (.A(clknet_1_1__leaf_net823),
    .Y(net1018));
 sky130_fd_sc_hd__inv_16 net999_11 (.A(clknet_1_0__leaf_net823),
    .Y(net1019));
 sky130_fd_sc_hd__inv_16 net999_12 (.A(clknet_1_0__leaf_net823),
    .Y(net1020));
 sky130_fd_sc_hd__inv_6 c232_14 (.A(clknet_1_0__leaf_net913),
    .Y(net1022));
 sky130_fd_sc_hd__inv_6 c232_15 (.A(clknet_1_0__leaf_net913),
    .Y(net1023));
 sky130_fd_sc_hd__inv_6 c232_16 (.A(clknet_1_0__leaf_net913),
    .Y(net1024));
 sky130_fd_sc_hd__inv_6 c232_17 (.A(clknet_1_0__leaf_net913),
    .Y(net1025));
 sky130_fd_sc_hd__inv_6 c232_18 (.A(clknet_1_1__leaf_net913),
    .Y(net1026));
 sky130_fd_sc_hd__inv_6 c232_19 (.A(clknet_1_0__leaf_net913),
    .Y(net1027));
 sky130_fd_sc_hd__inv_6 c250_21 (.A(clknet_1_1__leaf_net913),
    .Y(net1029));
 sky130_fd_sc_hd__inv_6 c250_22 (.A(clknet_1_1__leaf_net913),
    .Y(net1030));
 sky130_fd_sc_hd__inv_6 c250_23 (.A(clknet_1_1__leaf_net913),
    .Y(net1031));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net914 (.A(net914),
    .X(clknet_0_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net914 (.A(clknet_0_net914),
    .X(clknet_1_0__leaf_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net914 (.A(clknet_0_net914),
    .X(clknet_1_1__leaf_net914));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net548 (.A(net548),
    .X(clknet_0_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net548 (.A(clknet_0_net548),
    .X(clknet_1_0__leaf_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net548 (.A(clknet_0_net548),
    .X(clknet_1_1__leaf_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net666 (.A(net666),
    .X(clknet_0_net666));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net666 (.A(clknet_0_net666),
    .X(clknet_1_0__leaf_net666));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net666 (.A(clknet_0_net666),
    .X(clknet_1_1__leaf_net666));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net665 (.A(net665),
    .X(clknet_0_net665));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net665 (.A(clknet_0_net665),
    .X(clknet_1_0__leaf_net665));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net665 (.A(clknet_0_net665),
    .X(clknet_1_1__leaf_net665));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net894 (.A(net894),
    .X(clknet_0_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net724 (.A(net724),
    .X(clknet_0_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net724 (.A(clknet_0_net724),
    .X(clknet_1_0__leaf_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net724 (.A(clknet_0_net724),
    .X(clknet_1_1__leaf_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net715 (.A(net715),
    .X(clknet_0_net715));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net715 (.A(clknet_0_net715),
    .X(clknet_1_0__leaf_net715));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net715 (.A(clknet_0_net715),
    .X(clknet_1_1__leaf_net715));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net711 (.A(net711),
    .X(clknet_0_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net711 (.A(clknet_0_net711),
    .X(clknet_1_0__leaf_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net711 (.A(clknet_0_net711),
    .X(clknet_1_1__leaf_net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net655 (.A(net655),
    .X(clknet_0_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net657 (.A(net657),
    .X(clknet_0_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_0__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_1__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net912 (.A(net912),
    .X(clknet_0_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_0__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net912 (.A(clknet_0_net912),
    .X(clknet_1_1__leaf_net912));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net662 (.A(net662),
    .X(clknet_0_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net662 (.A(clknet_0_net662),
    .X(clknet_1_0__leaf_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net662 (.A(clknet_0_net662),
    .X(clknet_1_1__leaf_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net664 (.A(net664),
    .X(clknet_0_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_0__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_1__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net409 (.A(net409),
    .X(clknet_0_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_1__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net460 (.A(net460),
    .X(clknet_0_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_0__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net460 (.A(clknet_0_net460),
    .X(clknet_1_1__leaf_net460));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net467 (.A(net467),
    .X(clknet_0_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net467 (.A(clknet_0_net467),
    .X(clknet_1_0__leaf_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net467 (.A(clknet_0_net467),
    .X(clknet_1_1__leaf_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net466 (.A(net466),
    .X(clknet_0_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net466 (.A(clknet_0_net466),
    .X(clknet_1_0__leaf_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net466 (.A(clknet_0_net466),
    .X(clknet_1_1__leaf_net466));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net593 (.A(net593),
    .X(clknet_0_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net593 (.A(clknet_0_net593),
    .X(clknet_1_0__leaf_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net593 (.A(clknet_0_net593),
    .X(clknet_1_1__leaf_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net583 (.A(net583),
    .X(clknet_0_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net583 (.A(clknet_0_net583),
    .X(clknet_1_0__leaf_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net583 (.A(clknet_0_net583),
    .X(clknet_1_1__leaf_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net464 (.A(net464),
    .X(clknet_0_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net728 (.A(net728),
    .X(clknet_0_net728));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net728 (.A(clknet_0_net728),
    .X(clknet_1_0__leaf_net728));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net728 (.A(clknet_0_net728),
    .X(clknet_1_1__leaf_net728));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net581 (.A(net581),
    .X(clknet_0_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_0__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_1__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net957 (.A(net957),
    .X(clknet_0_net957));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net957 (.A(clknet_0_net957),
    .X(clknet_1_0__leaf_net957));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net957 (.A(clknet_0_net957),
    .X(clknet_1_1__leaf_net957));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net580 (.A(net580),
    .X(clknet_0_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_0__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_1__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net472 (.A(net472),
    .X(clknet_0_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_0__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_1__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net461 (.A(net461),
    .X(clknet_0_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net461 (.A(clknet_0_net461),
    .X(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net461 (.A(clknet_0_net461),
    .X(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net621 (.A(net621),
    .X(clknet_0_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net621 (.A(clknet_0_net621),
    .X(clknet_1_0__leaf_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net621 (.A(clknet_0_net621),
    .X(clknet_1_1__leaf_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net613 (.A(net613),
    .X(clknet_0_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net613 (.A(clknet_0_net613),
    .X(clknet_1_0__leaf_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net613 (.A(clknet_0_net613),
    .X(clknet_1_1__leaf_net613));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net611 (.A(net611),
    .X(clknet_0_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_0__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_1__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net486 (.A(net486),
    .X(clknet_0_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net486 (.A(clknet_0_net486),
    .X(clknet_1_0__leaf_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net486 (.A(clknet_0_net486),
    .X(clknet_1_1__leaf_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net459 (.A(net459),
    .X(clknet_0_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_0__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_1__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net822 (.A(net822),
    .X(clknet_0_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net822 (.A(clknet_0_net822),
    .X(clknet_1_0__leaf_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net822 (.A(clknet_0_net822),
    .X(clknet_1_1__leaf_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net427 (.A(net427),
    .X(clknet_0_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_0__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net427 (.A(clknet_0_net427),
    .X(clknet_1_1__leaf_net427));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net430 (.A(net430),
    .X(clknet_0_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net430 (.A(clknet_0_net430),
    .X(clknet_1_0__leaf_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net430 (.A(clknet_0_net430),
    .X(clknet_1_1__leaf_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net420 (.A(net420),
    .X(clknet_0_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_0__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net420 (.A(clknet_0_net420),
    .X(clknet_1_1__leaf_net420));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net554 (.A(net554),
    .X(clknet_0_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net554 (.A(net1039),
    .X(clknet_1_0__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_1__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net678 (.A(net678),
    .X(clknet_0_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net678 (.A(clknet_0_net678),
    .X(clknet_1_0__leaf_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net678 (.A(clknet_0_net678),
    .X(clknet_1_1__leaf_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net696 (.A(net696),
    .X(clknet_0_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net696 (.A(clknet_0_net696),
    .X(clknet_1_0__leaf_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net696 (.A(clknet_0_net696),
    .X(clknet_1_1__leaf_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net557 (.A(net557),
    .X(clknet_0_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_0__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_1__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net579 (.A(net579),
    .X(clknet_0_net579));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net579 (.A(clknet_0_net579),
    .X(clknet_1_0__leaf_net579));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net579 (.A(clknet_0_net579),
    .X(clknet_1_1__leaf_net579));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net913 (.A(net913),
    .X(clknet_0_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net913 (.A(clknet_0_net913),
    .X(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net913 (.A(clknet_0_net913),
    .X(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net234 (.A(net234),
    .X(clknet_0_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net240 (.A(net240),
    .X(clknet_0_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net240 (.A(clknet_0_net240),
    .X(clknet_1_0__leaf_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net240 (.A(clknet_0_net240),
    .X(clknet_1_1__leaf_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net841 (.A(net841),
    .X(clknet_0_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net841 (.A(clknet_0_net841),
    .X(clknet_1_0__leaf_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net841 (.A(clknet_0_net841),
    .X(clknet_1_1__leaf_net841));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net499 (.A(net499),
    .X(clknet_0_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_0__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_1__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net502 (.A(net502),
    .X(clknet_0_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_0__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_1__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net875 (.A(net875),
    .X(clknet_0_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net875 (.A(clknet_0_net875),
    .X(clknet_1_0__leaf_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net875 (.A(clknet_0_net875),
    .X(clknet_1_1__leaf_net875));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net214 (.A(net214),
    .X(clknet_0_net214));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net214 (.A(clknet_0_net214),
    .X(clknet_1_0__leaf_net214));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net214 (.A(clknet_0_net214),
    .X(clknet_1_1__leaf_net214));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net858 (.A(net858),
    .X(clknet_0_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net858 (.A(clknet_0_net858),
    .X(clknet_1_0__leaf_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net858 (.A(clknet_0_net858),
    .X(clknet_1_1__leaf_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net223 (.A(net223),
    .X(clknet_0_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_0__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_1__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net241 (.A(net241),
    .X(clknet_0_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_0__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_1__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net839 (.A(net839),
    .X(clknet_0_net839));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net839 (.A(clknet_0_net839),
    .X(clknet_1_0__leaf_net839));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net839 (.A(clknet_0_net839),
    .X(clknet_1_1__leaf_net839));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net222 (.A(net222),
    .X(clknet_0_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_0__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_1__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net352 (.A(net352),
    .X(clknet_0_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net892 (.A(net892),
    .X(clknet_0_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_0__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_1__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net876 (.A(net876),
    .X(clknet_0_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net876 (.A(clknet_0_net876),
    .X(clknet_1_0__leaf_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net876 (.A(clknet_0_net876),
    .X(clknet_1_1__leaf_net876));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net534 (.A(net534),
    .X(clknet_0_net534));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net534 (.A(clknet_0_net534),
    .X(clknet_1_0__leaf_net534));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net534 (.A(clknet_0_net534),
    .X(clknet_1_1__leaf_net534));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net645 (.A(net645),
    .X(clknet_0_net645));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net645 (.A(clknet_0_net645),
    .X(clknet_1_0__leaf_net645));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net645 (.A(clknet_0_net645),
    .X(clknet_1_1__leaf_net645));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net629 (.A(net629),
    .X(clknet_0_net629));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net629 (.A(clknet_0_net629),
    .X(clknet_1_0__leaf_net629));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net629 (.A(clknet_0_net629),
    .X(clknet_1_1__leaf_net629));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net639 (.A(net639),
    .X(clknet_0_net639));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net639 (.A(clknet_0_net639),
    .X(clknet_1_0__leaf_net639));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net639 (.A(clknet_0_net639),
    .X(clknet_1_1__leaf_net639));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net641 (.A(net641),
    .X(clknet_0_net641));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net641 (.A(clknet_0_net641),
    .X(clknet_1_0__leaf_net641));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net641 (.A(clknet_0_net641),
    .X(clknet_1_1__leaf_net641));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net533 (.A(net533),
    .X(clknet_0_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net533 (.A(clknet_0_net533),
    .X(clknet_1_0__leaf_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net533 (.A(clknet_0_net533),
    .X(clknet_1_1__leaf_net533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net556 (.A(net556),
    .X(clknet_0_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_0__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_1__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net649 (.A(net649),
    .X(clknet_0_net649));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net649 (.A(clknet_0_net649),
    .X(clknet_1_0__leaf_net649));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net649 (.A(clknet_0_net649),
    .X(clknet_1_1__leaf_net649));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net540 (.A(net540),
    .X(clknet_0_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_0__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_1__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net532 (.A(net532),
    .X(clknet_0_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_0__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_1__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net967 (.A(net967),
    .X(clknet_0_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net967 (.A(clknet_0_net967),
    .X(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net967 (.A(clknet_0_net967),
    .X(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net679 (.A(net679),
    .X(clknet_0_net679));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net679 (.A(clknet_0_net679),
    .X(clknet_1_0__leaf_net679));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net679 (.A(clknet_0_net679),
    .X(clknet_1_1__leaf_net679));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net674 (.A(net674),
    .X(clknet_0_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net674 (.A(clknet_0_net674),
    .X(clknet_1_0__leaf_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net674 (.A(clknet_0_net674),
    .X(clknet_1_1__leaf_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net574 (.A(net574),
    .X(clknet_0_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_0__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_1__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net578 (.A(net578),
    .X(clknet_0_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net578 (.A(clknet_0_net578),
    .X(clknet_1_0__leaf_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net578 (.A(clknet_0_net578),
    .X(clknet_1_1__leaf_net578));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net821 (.A(net821),
    .X(clknet_0_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net821 (.A(clknet_0_net821),
    .X(clknet_1_0__leaf_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net821 (.A(clknet_0_net821),
    .X(clknet_1_1__leaf_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net440 (.A(net440),
    .X(clknet_0_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_0__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_1__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net441 (.A(net441),
    .X(clknet_0_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net441 (.A(clknet_0_net441),
    .X(clknet_1_0__leaf_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net441 (.A(clknet_0_net441),
    .X(clknet_1_1__leaf_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net584 (.A(net584),
    .X(clknet_0_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_0__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net972 (.A(net972),
    .X(clknet_0_net972));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net972 (.A(clknet_0_net972),
    .X(clknet_1_0__leaf_net972));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net972 (.A(clknet_0_net972),
    .X(clknet_1_1__leaf_net972));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net840 (.A(net840),
    .X(clknet_0_net840));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net840 (.A(clknet_0_net840),
    .X(clknet_1_0__leaf_net840));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net840 (.A(clknet_0_net840),
    .X(clknet_1_1__leaf_net840));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net823 (.A(net823),
    .X(clknet_0_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net83 (.A(net83),
    .X(clknet_0_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net83 (.A(clknet_0_net83),
    .X(clknet_1_0__leaf_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net83 (.A(clknet_0_net83),
    .X(clknet_1_1__leaf_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net85 (.A(net85),
    .X(clknet_0_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net85 (.A(clknet_0_net85),
    .X(clknet_1_0__leaf_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net85 (.A(clknet_0_net85),
    .X(clknet_1_1__leaf_net85));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net103 (.A(net103),
    .X(clknet_0_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net103 (.A(clknet_0_net103),
    .X(clknet_1_0__leaf_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net103 (.A(clknet_0_net103),
    .X(clknet_1_1__leaf_net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net365 (.A(net365),
    .X(clknet_0_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net370 (.A(net370),
    .X(clknet_0_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_0__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net367 (.A(net367),
    .X(clknet_0_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_0__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_1__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net81 (.A(net81),
    .X(clknet_0_net81));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net81 (.A(clknet_0_net81),
    .X(clknet_1_0__leaf_net81));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net81 (.A(clknet_0_net81),
    .X(clknet_1_1__leaf_net81));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net339 (.A(net339),
    .X(clknet_0_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net339 (.A(clknet_0_net339),
    .X(clknet_1_0__leaf_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net339 (.A(clknet_0_net339),
    .X(clknet_1_1__leaf_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net210 (.A(net210),
    .X(clknet_0_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_0__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net210 (.A(clknet_0_net210),
    .X(clknet_1_1__leaf_net210));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net78 (.A(net78),
    .X(clknet_0_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net78 (.A(clknet_0_net78),
    .X(clknet_1_0__leaf_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net78 (.A(clknet_0_net78),
    .X(clknet_1_1__leaf_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net346 (.A(net346),
    .X(clknet_0_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net478 (.A(net478),
    .X(clknet_0_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_0__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_1__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net201 (.A(net201),
    .X(clknet_0_net201));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net201 (.A(clknet_0_net201),
    .X(clknet_1_0__leaf_net201));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net201 (.A(clknet_0_net201),
    .X(clknet_1_1__leaf_net201));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net471 (.A(net471),
    .X(clknet_0_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_0__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_1__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net89 (.A(net89),
    .X(clknet_0_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net89 (.A(clknet_0_net89),
    .X(clknet_1_0__leaf_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net89 (.A(clknet_0_net89),
    .X(clknet_1_1__leaf_net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net364 (.A(net364),
    .X(clknet_0_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net364 (.A(clknet_0_net364),
    .X(clknet_1_0__leaf_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net364 (.A(clknet_0_net364),
    .X(clknet_1_1__leaf_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net501 (.A(net501),
    .X(clknet_0_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_0__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_1__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net225 (.A(net225),
    .X(clknet_0_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net225 (.A(clknet_0_net225),
    .X(clknet_1_0__leaf_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net225 (.A(clknet_0_net225),
    .X(clknet_1_1__leaf_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net227 (.A(net227),
    .X(clknet_0_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net227 (.A(clknet_0_net227),
    .X(clknet_1_0__leaf_net227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net227 (.A(clknet_0_net227),
    .X(clknet_1_1__leaf_net227));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer1 (.A(net1065),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1065),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net231),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net121),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net124),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net970),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net1008),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer8 (.A(net1035),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer9 (.A(net1036),
    .X(net1037));
 sky130_fd_sc_hd__clkbuf_1 clone10 (.A(net1007),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(clknet_0_net554),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net1003),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net952),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net653),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net485),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net319),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net811),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net871),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net693),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net961),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net796),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net87),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net955),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net350),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net306),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net940),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net864),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net850),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net96),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net949),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net488),
    .X(net1059));
 sky130_fd_sc_hd__clkbuf_1 wire1 (.A(net770),
    .X(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_S0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A3 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_C_N (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_S0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_SCE (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_C (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_Y (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A3 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_RESET_B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_D_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_Y (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_D1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B_N (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_C (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_Y (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A_N (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B_N (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_C_N (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_D1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_D (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_C1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_C_N (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B_N (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_Y (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A_N (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_SET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_SCE (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_D (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_C_N (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_Y (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_SCE (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_C_N (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_C (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_Y (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_C (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_Y (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A3 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A3 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A_N (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_SCE (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_D (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_RESET_B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_D (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_Q (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_C_N (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_X (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A0 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A3 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A_N (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_Q (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B_N (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_Y (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_Y (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_RESET_B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_Y (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_D (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B_N (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_SCD (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_D1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_SCE (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SCD (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_D1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_D1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A3 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_D_N (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_D1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_Y (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_X (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_C1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_C_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_Y (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_Y (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_SCD (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S0 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S0 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_D (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_D (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_SCD (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_C_N (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A_N (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_X (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A3 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_C_N (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A_N (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_Y (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A0 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_C (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_C1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B_N (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_C_N (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_SCE (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_S0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_SCD (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_C_N (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_SCD (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_SCE (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_D (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_SET_B (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_RESET_B (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_X (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B_N (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A3 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_Y (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_C_N (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_D1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_RESET_B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_D_N (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S0 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_C1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_Q_N (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_C1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_Q (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_C1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_Q_N (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_RESET_B (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B_N (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_Q (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_RESET_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_X (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold16_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_D1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_SCD (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_Y (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A3 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_SCD (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_D (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_Y (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_S1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_Q_N (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_C_N (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_D (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_X (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A3 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A0 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A3 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_X (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_RESET_B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_A1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A3 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_X (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_RESET_B (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Y (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_RESET_B (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_B (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_X (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A_N (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_Y (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_SCD (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_Y (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_B (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A_N (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_C1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_C (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_DE (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_C (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_Y (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_RESET_B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_C_N (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_D (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_D1 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_D_N (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_C (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_Y (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_A1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_SET_B (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A_N (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_C_N (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B_N (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_Y (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_Y (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_D (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_SCD (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_RESET_B (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_X (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_B1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_C_N (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_Q (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_DE (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_Y (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A0 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_C1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_X (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_C1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_D (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_C1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_D_N (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_SET_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_C_N (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B_N (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_Y (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_C1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap76_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_Y (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_C_N (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_C1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_Y (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_B1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_C1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SCD (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_C_N (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_Y (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_Y (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_C_N (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_B (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_C1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_SCD (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B_N (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A_N (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_X (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_D1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_B_N (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_SCD (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_Q_N (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A_N (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_Q (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_SET_B (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_RESET_B (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_D (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_X (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_SCE (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_D (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S0 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_X (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A2 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_C_N (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_D_N (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_X (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_SCE (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_D (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_D_N (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_Y (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_Y (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_SET_B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_Y (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_SCE (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_X (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_SET_B (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_B (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_SCE (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_Q (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_X (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net578_A (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_X (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_C (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_RESET_B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_D (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A3 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_C (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_Y (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A3 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_S1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_D (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_SCE (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_C1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_D1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_Y (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A0 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_RESET_B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_X (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_C_N (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_D (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_X (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net665_A (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_X (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_B1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_Q (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_Q (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_Y (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_RESET_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_Y (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold17_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_Q (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_C (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_SCE (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net823_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_GCLK (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_Q (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_s847_Q (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_Q_N (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_Q (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_S1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_C_N (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_D1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_Q_N (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_S1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_C (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_C_N (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_Q (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_SCE (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_D_N (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_D1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_Q (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_SET_B (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_Q (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_Q (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_D1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_D1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_D_N (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_Q_N (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_Q (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_C (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_D (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_S0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_S1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_C1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_C (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A_N (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B_N (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_D1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_C1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_C (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B_N (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_SET_B (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_SCE (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_SCE (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_C_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_A_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_B (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_B1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_A0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_SCE (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_D (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_C_N (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold26_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A_N (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_B_N (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_C1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_D_N (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B_N (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_D_N (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_SCE (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold30_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_Q (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold13_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold20_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_Q (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_D1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_SET_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_D1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_D1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_B1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_RESET_B (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_Q (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net967_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_GCLK (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_D1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_Y (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_C (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_Q (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net972_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_GCLK (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire52_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_SCE (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_SCE (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_C_N (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_SCD (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_SCE (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_S1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_SCD (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_SCE (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_B (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_SET_B (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_RESET_B (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_SCE (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_C_N (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_C_N (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_D1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_D_N (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SCE (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_C_N (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_SCD (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_D1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_C_N (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_C (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_D1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_C_N (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_D_N (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_C (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_C (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_C1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_SCE (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_SET_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_C (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_D_N (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_SCD (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap62_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_B1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_B (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_C (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_C (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_D1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_C1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_B1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_C_N (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A3 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A3 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_C1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SCE (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_SET_B (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_RESET_B (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_C_N (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap67_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire69_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap67_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap68_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap71_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap70_A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire73_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire72_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap74_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_C_N (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_SCE (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_SCD (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_C (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_SCE (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_C1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_D_N (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_D_N (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap76_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_D1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_B_N (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_D_N (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_D_N (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_SCE (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_C_N (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_D_N (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_SCD (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_D_N (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_SCD (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_C_N (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_S0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_D1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_D_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_C_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_C_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_D_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_SET_B (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_SET_B (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_C (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_D1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_C_N (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_D_N (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_D_N (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold12_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_C1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_D_N (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_SCE (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_A (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_SCE (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_SCD (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_D_N (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_B (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_C (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_D_N (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s846_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s847_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s843_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s848_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s844_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s845_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s850_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s851_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_SLEEP_B (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_SCD (.DIODE(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net461_X (.DIODE(clknet_1_0__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_C1 (.DIODE(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_B1 (.DIODE(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_B1 (.DIODE(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_C1 (.DIODE(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net461_X (.DIODE(clknet_1_1__leaf_net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(clknet_1_0__leaf_net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_S0 (.DIODE(clknet_1_0__leaf_net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net822_X (.DIODE(clknet_1_0__leaf_net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net967_A (.DIODE(clknet_0_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net967_A (.DIODE(clknet_0_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net967_X (.DIODE(clknet_0_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B (.DIODE(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SET_B (.DIODE(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_C (.DIODE(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_S1 (.DIODE(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net967_X (.DIODE(clknet_1_0__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_S1 (.DIODE(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_S1 (.DIODE(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_D1 (.DIODE(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net967_X (.DIODE(clknet_1_1__leaf_net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_C_N (.DIODE(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_B (.DIODE(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_B (.DIODE(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_C1 (.DIODE(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net562_X (.DIODE(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net972_A (.DIODE(clknet_0_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net972_A (.DIODE(clknet_0_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net972_X (.DIODE(clknet_0_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S1 (.DIODE(clknet_1_0__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_C (.DIODE(clknet_1_0__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_D1 (.DIODE(clknet_1_0__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_SET_B (.DIODE(clknet_1_0__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net972_X (.DIODE(clknet_1_0__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_D1 (.DIODE(clknet_1_1__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_S1 (.DIODE(clknet_1_1__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(clknet_1_1__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_D1 (.DIODE(clknet_1_1__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(clknet_1_1__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net972_X (.DIODE(clknet_1_1__leaf_net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net823_A (.DIODE(clknet_0_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net823_A (.DIODE(clknet_0_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net823_X (.DIODE(clknet_0_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_B (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_1_A (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_7_A (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_8_A (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_9_A (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_11_A (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_12_A (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net823_X (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_2_A (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_3_A (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_4_A (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_5_A (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_6_A (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_10_A (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net823_X (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_D_N (.DIODE(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_B1 (.DIODE(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net346_X (.DIODE(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(clknet_1_0__leaf_net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(clknet_1_0__leaf_net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B (.DIODE(clknet_1_0__leaf_net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_D_N (.DIODE(clknet_1_0__leaf_net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net201_X (.DIODE(clknet_1_0__leaf_net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(clknet_1_1__leaf_net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A2 (.DIODE(clknet_1_1__leaf_net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A0 (.DIODE(clknet_1_1__leaf_net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A0 (.DIODE(clknet_1_1__leaf_net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net201_X (.DIODE(clknet_1_1__leaf_net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A2 (.DIODE(clknet_1_0__leaf_net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A2 (.DIODE(clknet_1_0__leaf_net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A3 (.DIODE(clknet_1_0__leaf_net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A2 (.DIODE(clknet_1_0__leaf_net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A2 (.DIODE(clknet_1_0__leaf_net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net364_X (.DIODE(clknet_1_0__leaf_net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_B (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_D1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_C1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_RESET_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_A (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold26_X (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net112));
 sky130_fd_sc_hd__and2_1 clone1 (.A(net1063),
    .B(net245),
    .X(net1061));
 sky130_fd_sc_hd__and2_1 clone2 (.A(net1063),
    .B(net245),
    .X(net1062));
 sky130_fd_sc_hd__and2b_1 clone3 (.A_N(net944),
    .B(net995),
    .X(net1063));
 sky130_fd_sc_hd__clkbuf_1 clone4 (.A(net1008),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net121),
    .X(net1065));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
