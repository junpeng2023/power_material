module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net1003;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net1008;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net1010;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire clknet_0_clk;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net1013;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1009;
 wire net1011;
 wire net1012;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net920;
 wire clknet_1_0__leaf_net920;
 wire clknet_1_1__leaf_net920;
 wire clknet_0_net655;
 wire clknet_1_0__leaf_net655;
 wire clknet_1_1__leaf_net655;
 wire clknet_0_net673;
 wire clknet_1_0__leaf_net673;
 wire clknet_1_1__leaf_net673;
 wire clknet_0_net677;
 wire clknet_1_0__leaf_net677;
 wire clknet_1_1__leaf_net677;
 wire clknet_0_net756;
 wire clknet_1_0__leaf_net756;
 wire clknet_1_1__leaf_net756;
 wire clknet_0_net630;
 wire clknet_1_0__leaf_net630;
 wire clknet_1_1__leaf_net630;
 wire clknet_0_net634;
 wire clknet_1_0__leaf_net634;
 wire clknet_1_1__leaf_net634;
 wire clknet_0_net640;
 wire clknet_1_0__leaf_net640;
 wire clknet_1_1__leaf_net640;
 wire clknet_0_net622;
 wire clknet_1_0__leaf_net622;
 wire clknet_1_1__leaf_net622;
 wire clknet_0_net919;
 wire clknet_1_0__leaf_net919;
 wire clknet_1_1__leaf_net919;
 wire clknet_0_net631;
 wire clknet_1_0__leaf_net631;
 wire clknet_1_1__leaf_net631;
 wire clknet_0_net544;
 wire clknet_1_0__leaf_net544;
 wire clknet_1_1__leaf_net544;
 wire clknet_0_net324;
 wire clknet_1_0__leaf_net324;
 wire clknet_1_1__leaf_net324;
 wire clknet_0_net475;
 wire clknet_1_0__leaf_net475;
 wire clknet_1_1__leaf_net475;
 wire clknet_0_net843;
 wire clknet_1_0__leaf_net843;
 wire clknet_1_1__leaf_net843;
 wire clknet_0_net472;
 wire clknet_1_0__leaf_net472;
 wire clknet_1_1__leaf_net472;
 wire clknet_0_net956;
 wire clknet_1_0__leaf_net956;
 wire clknet_1_1__leaf_net956;
 wire clknet_0_net478;
 wire clknet_1_0__leaf_net478;
 wire clknet_1_1__leaf_net478;
 wire clknet_0_net476;
 wire clknet_1_0__leaf_net476;
 wire clknet_1_1__leaf_net476;
 wire clknet_0_net327;
 wire clknet_1_0__leaf_net327;
 wire clknet_1_1__leaf_net327;
 wire clknet_0_net531;
 wire clknet_1_0__leaf_net531;
 wire clknet_1_1__leaf_net531;
 wire clknet_0_net553;
 wire clknet_1_0__leaf_net553;
 wire clknet_1_1__leaf_net553;
 wire clknet_0_net603;
 wire clknet_1_0__leaf_net603;
 wire clknet_1_1__leaf_net603;
 wire clknet_0_net951;
 wire clknet_1_0__leaf_net951;
 wire clknet_1_1__leaf_net951;
 wire clknet_0_net612;
 wire clknet_1_0__leaf_net612;
 wire clknet_1_1__leaf_net612;
 wire clknet_0_net947;
 wire clknet_1_0__leaf_net947;
 wire clknet_1_1__leaf_net947;
 wire clknet_0_net608;
 wire clknet_1_0__leaf_net608;
 wire clknet_1_1__leaf_net608;
 wire clknet_0_net605;
 wire clknet_1_0__leaf_net605;
 wire clknet_1_1__leaf_net605;
 wire clknet_0_net609;
 wire clknet_1_0__leaf_net609;
 wire clknet_1_1__leaf_net609;
 wire clknet_0_net602;
 wire clknet_1_0__leaf_net602;
 wire clknet_1_1__leaf_net602;
 wire clknet_0_net388;
 wire clknet_1_0__leaf_net388;
 wire clknet_1_1__leaf_net388;
 wire clknet_0_net508;
 wire clknet_1_0__leaf_net508;
 wire clknet_1_1__leaf_net508;
 wire clknet_0_net519;
 wire clknet_1_0__leaf_net519;
 wire clknet_1_1__leaf_net519;
 wire clknet_0_net513;
 wire clknet_1_0__leaf_net513;
 wire clknet_1_1__leaf_net513;
 wire clknet_0_net664;
 wire clknet_1_0__leaf_net664;
 wire clknet_1_1__leaf_net664;
 wire clknet_0_net621;
 wire clknet_1_0__leaf_net621;
 wire clknet_1_1__leaf_net621;
 wire clknet_0_net565;
 wire clknet_1_0__leaf_net565;
 wire clknet_1_1__leaf_net565;
 wire clknet_0_net808;
 wire clknet_1_0__leaf_net808;
 wire clknet_1_1__leaf_net808;
 wire clknet_0_net562;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_1__leaf_net562;
 wire clknet_0_net529;
 wire clknet_1_0__leaf_net529;
 wire clknet_1_1__leaf_net529;
 wire clknet_0_net862;
 wire clknet_1_0__leaf_net862;
 wire clknet_1_1__leaf_net862;
 wire clknet_0_net638;
 wire clknet_1_0__leaf_net638;
 wire clknet_1_1__leaf_net638;
 wire clknet_0_net637;
 wire clknet_1_0__leaf_net637;
 wire clknet_1_1__leaf_net637;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net390;
 wire clknet_1_0__leaf_net390;
 wire clknet_1_1__leaf_net390;
 wire clknet_0_net898;
 wire clknet_1_0__leaf_net898;
 wire clknet_1_1__leaf_net898;
 wire clknet_0_net168;
 wire clknet_1_0__leaf_net168;
 wire clknet_1_1__leaf_net168;
 wire clknet_0_net223;
 wire clknet_1_0__leaf_net223;
 wire clknet_1_1__leaf_net223;
 wire clknet_0_net238;
 wire clknet_1_0__leaf_net238;
 wire clknet_1_1__leaf_net238;
 wire clknet_0_net950;
 wire clknet_1_0__leaf_net950;
 wire clknet_1_1__leaf_net950;
 wire clknet_0_net970;
 wire clknet_1_0__leaf_net970;
 wire clknet_1_1__leaf_net970;
 wire clknet_0_net806;
 wire clknet_1_0__leaf_net806;
 wire clknet_1_1__leaf_net806;
 wire clknet_0_net233;
 wire clknet_1_0__leaf_net233;
 wire clknet_1_1__leaf_net233;
 wire clknet_0_net165;
 wire clknet_1_0__leaf_net165;
 wire clknet_1_1__leaf_net165;
 wire clknet_0_net422;
 wire clknet_1_0__leaf_net422;
 wire clknet_1_1__leaf_net422;
 wire clknet_0_net426;
 wire clknet_1_0__leaf_net426;
 wire clknet_1_1__leaf_net426;
 wire clknet_0_net558;
 wire clknet_1_0__leaf_net558;
 wire clknet_1_1__leaf_net558;
 wire clknet_0_net550;
 wire clknet_1_0__leaf_net550;
 wire clknet_1_1__leaf_net550;
 wire clknet_0_net659;
 wire clknet_1_0__leaf_net659;
 wire clknet_1_1__leaf_net659;
 wire clknet_0_net702;
 wire clknet_1_0__leaf_net702;
 wire clknet_1_1__leaf_net702;
 wire clknet_0_net547;
 wire clknet_1_0__leaf_net547;
 wire clknet_1_1__leaf_net547;
 wire clknet_0_net549;
 wire clknet_1_0__leaf_net549;
 wire clknet_1_1__leaf_net549;
 wire clknet_0_net860;
 wire clknet_1_0__leaf_net860;
 wire clknet_1_1__leaf_net860;
 wire clknet_0_net428;
 wire clknet_1_0__leaf_net428;
 wire clknet_1_1__leaf_net428;
 wire clknet_0_net430;
 wire clknet_1_0__leaf_net430;
 wire clknet_1_1__leaf_net430;
 wire clknet_0_net295;
 wire clknet_1_0__leaf_net295;
 wire clknet_1_1__leaf_net295;
 wire clknet_0_net313;
 wire clknet_1_0__leaf_net313;
 wire clknet_1_1__leaf_net313;
 wire clknet_0_net171;
 wire clknet_1_0__leaf_net171;
 wire clknet_1_1__leaf_net171;
 wire clknet_0_net585;
 wire clknet_1_0__leaf_net585;
 wire clknet_1_1__leaf_net585;
 wire clknet_0_net587;
 wire clknet_1_0__leaf_net587;
 wire clknet_1_1__leaf_net587;
 wire clknet_0_net576;
 wire clknet_1_0__leaf_net576;
 wire clknet_1_1__leaf_net576;
 wire clknet_0_net589;
 wire clknet_1_0__leaf_net589;
 wire clknet_1_1__leaf_net589;
 wire clknet_0_net167;
 wire clknet_1_0__leaf_net167;
 wire clknet_1_1__leaf_net167;
 wire clknet_0_net435;
 wire clknet_1_0__leaf_net435;
 wire clknet_1_1__leaf_net435;
 wire clknet_0_net561;
 wire clknet_1_0__leaf_net561;
 wire clknet_1_1__leaf_net561;
 wire clknet_0_net557;
 wire clknet_1_0__leaf_net557;
 wire clknet_1_1__leaf_net557;
 wire clknet_0_net170;
 wire clknet_1_0__leaf_net170;
 wire clknet_1_1__leaf_net170;
 wire clknet_0_net205;
 wire clknet_1_0__leaf_net205;
 wire clknet_1_1__leaf_net205;
 wire clknet_0_net331;
 wire clknet_1_0__leaf_net331;
 wire clknet_1_1__leaf_net331;
 wire clknet_0_net823;
 wire clknet_1_0__leaf_net823;
 wire clknet_1_1__leaf_net823;
 wire clknet_0_net463;
 wire clknet_1_0__leaf_net463;
 wire clknet_1_1__leaf_net463;
 wire clknet_0_net596;
 wire clknet_1_0__leaf_net596;
 wire clknet_1_1__leaf_net596;
 wire clknet_0_net824;
 wire clknet_1_0__leaf_net824;
 wire clknet_1_1__leaf_net824;
 wire clknet_0_net369;
 wire clknet_1_0__leaf_net369;
 wire clknet_1_1__leaf_net369;
 wire clknet_0_net358;
 wire clknet_1_0__leaf_net358;
 wire clknet_1_1__leaf_net358;
 wire clknet_0_net966;
 wire clknet_1_0__leaf_net966;
 wire clknet_1_1__leaf_net966;
 wire clknet_0_net958;
 wire clknet_1_0__leaf_net958;
 wire clknet_1_1__leaf_net958;
 wire clknet_0_net594;
 wire clknet_1_0__leaf_net594;
 wire clknet_1_1__leaf_net594;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net341;
 wire clknet_1_0__leaf_net341;
 wire clknet_1_1__leaf_net341;
 wire clknet_0_net207;
 wire clknet_1_0__leaf_net207;
 wire clknet_1_1__leaf_net207;
 wire clknet_0_net211;
 wire clknet_1_0__leaf_net211;
 wire clknet_1_1__leaf_net211;
 wire clknet_0_net844;
 wire clknet_1_0__leaf_net844;
 wire clknet_1_1__leaf_net844;
 wire clknet_0_net198;
 wire clknet_1_0__leaf_net198;
 wire clknet_1_1__leaf_net198;
 wire clknet_0_net202;
 wire clknet_1_0__leaf_net202;
 wire clknet_1_1__leaf_net202;
 wire clknet_0_net213;
 wire clknet_1_0__leaf_net213;
 wire clknet_1_1__leaf_net213;
 wire clknet_0_net208;
 wire clknet_1_0__leaf_net208;
 wire clknet_1_1__leaf_net208;
 wire clknet_0_net897;
 wire clknet_1_0__leaf_net897;
 wire clknet_1_1__leaf_net897;
 wire clknet_0_net398;
 wire clknet_1_0__leaf_net398;
 wire clknet_1_1__leaf_net398;
 wire clknet_0_net446;
 wire clknet_1_0__leaf_net446;
 wire clknet_1_1__leaf_net446;
 wire clknet_0_net694;
 wire clknet_1_0__leaf_net694;
 wire clknet_1_1__leaf_net694;
 wire clknet_0_net718;
 wire clknet_1_0__leaf_net718;
 wire clknet_1_1__leaf_net718;
 wire clknet_0_net593;
 wire clknet_1_0__leaf_net593;
 wire clknet_1_1__leaf_net593;
 wire clknet_0_net842;
 wire clknet_1_0__leaf_net842;
 wire clknet_1_1__leaf_net842;
 wire clknet_0_net586;
 wire clknet_1_0__leaf_net586;
 wire clknet_1_1__leaf_net586;
 wire clknet_0_net405;
 wire clknet_1_0__leaf_net405;
 wire clknet_1_1__leaf_net405;
 wire clknet_0_net395;
 wire clknet_1_0__leaf_net395;
 wire clknet_1_1__leaf_net395;
 wire clknet_0_net416;
 wire clknet_1_0__leaf_net416;
 wire clknet_1_1__leaf_net416;
 wire clknet_0_net431;
 wire clknet_1_0__leaf_net431;
 wire clknet_1_1__leaf_net431;
 wire clknet_0_net425;
 wire clknet_1_0__leaf_net425;
 wire clknet_1_1__leaf_net425;
 wire clknet_0_net432;
 wire clknet_1_0__leaf_net432;
 wire clknet_1_1__leaf_net432;
 wire clknet_0_net861;
 wire clknet_1_0__leaf_net861;
 wire clknet_1_1__leaf_net861;
 wire net154;
 wire net162;
 wire net323;
 wire net625;
 wire net635;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;

 sky130_fd_sc_hd__nand2b_1 c100 (.A_N(net69),
    .B(net63),
    .Y(net74));
 sky130_fd_sc_hd__and2b_1 c101 (.A_N(net42),
    .B(net74),
    .X(net75));
 sky130_fd_sc_hd__or2_4 c102 (.A(net74),
    .B(net68),
    .X(net76));
 sky130_fd_sc_hd__and2b_1 c103 (.A_N(net67),
    .B(net74),
    .X(net77));
 sky130_fd_sc_hd__or2_1 c104 (.A(net941),
    .B(net17),
    .X(net78));
 sky130_fd_sc_hd__nor2b_4 c105 (.A(net928),
    .B_N(net68),
    .Y(net79));
 sky130_fd_sc_hd__nand2_1 c106 (.A(net68),
    .B(net79),
    .Y(net80));
 sky130_fd_sc_hd__nand2_1 c107 (.A(net72),
    .B(net75),
    .Y(net81));
 sky130_fd_sc_hd__or2b_2 c108 (.A(net73),
    .B_N(net75),
    .X(net82));
 sky130_fd_sc_hd__and3_2 c109 (.A(net80),
    .B(net81),
    .C(net62),
    .X(net83));
 sky130_fd_sc_hd__nand2b_1 c110 (.A_N(net70),
    .B(net63),
    .Y(net84));
 sky130_fd_sc_hd__or2_4 c111 (.A(net926),
    .B(net82),
    .X(net85));
 sky130_fd_sc_hd__inv_1 c112 (.A(net732),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 c113 (.A(net912),
    .Y(net87));
 sky130_fd_sc_hd__and2b_4 c114 (.A_N(net86),
    .B(net84),
    .X(net955));
 sky130_fd_sc_hd__nand2_1 c115 (.A(net33),
    .B(net86),
    .Y(net88));
 sky130_fd_sc_hd__or2b_1 c116 (.A(net35),
    .B_N(net85),
    .X(net89));
 sky130_fd_sc_hd__or2b_1 c117 (.A(net17),
    .B_N(net85),
    .X(net90));
 sky130_fd_sc_hd__nand2b_1 c118 (.A_N(net58),
    .B(net64),
    .Y(net91));
 sky130_fd_sc_hd__inv_4 c119 (.A(net732),
    .Y(net92));
 sky130_fd_sc_hd__inv_6 c120 (.A(net1018),
    .Y(net93));
 sky130_fd_sc_hd__inv_12 c121 (.A(net814),
    .Y(net94));
 sky130_fd_sc_hd__or2_1 c122 (.A(net87),
    .B(net63),
    .X(net95));
 sky130_fd_sc_hd__or2_1 c123 (.A(net85),
    .B(net798),
    .X(net96));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net84),
    .A1(net30),
    .A2(net92),
    .A3(net58),
    .S0(net32),
    .S1(net955),
    .X(net97));
 sky130_fd_sc_hd__nor3b_1 c125 (.A(net35),
    .B(net94),
    .C_N(net787),
    .Y(net98));
 sky130_fd_sc_hd__nand2b_1 c126 (.A_N(net69),
    .B(net93),
    .Y(net99));
 sky130_fd_sc_hd__inv_2 c127 (.A(net911),
    .Y(net100));
 sky130_fd_sc_hd__clkbuf_2 c128 (.A(net918),
    .X(net101));
 sky130_fd_sc_hd__mux4_2 c129 (.A0(net99),
    .A1(net98),
    .A2(net64),
    .A3(net101),
    .S0(net17),
    .S1(net162),
    .X(net102));
 sky130_fd_sc_hd__mux4_2 c130 (.A0(net93),
    .A1(net99),
    .A2(net94),
    .A3(net89),
    .S0(net101),
    .S1(net817),
    .X(net103));
 sky130_fd_sc_hd__mux4_4 c131 (.A0(net89),
    .A1(net100),
    .A2(net101),
    .A3(net33),
    .S0(net85),
    .S1(net1030),
    .X(net104));
 sky130_fd_sc_hd__and2b_4 c132 (.A_N(net924),
    .B(net943),
    .X(net105));
 sky130_fd_sc_hd__nor2_2 c133 (.A(net944),
    .B(net932),
    .Y(net106));
 sky130_fd_sc_hd__or2_4 c134 (.A(net942),
    .B(net1000),
    .X(net107));
 sky130_fd_sc_hd__nor2b_2 c135 (.A(net931),
    .B_N(net927),
    .Y(net108));
 sky130_fd_sc_hd__nor2_2 c136 (.A(net929),
    .B(net1000),
    .Y(net109));
 sky130_fd_sc_hd__or2_1 c137 (.A(net922),
    .B(net929),
    .X(net110));
 sky130_fd_sc_hd__and2_2 c138 (.A(net108),
    .B(net930),
    .X(net111));
 sky130_fd_sc_hd__nand2_2 c139 (.A(net106),
    .B(net924),
    .Y(net112));
 sky130_fd_sc_hd__nand2_4 c140 (.A(net108),
    .B(net932),
    .Y(net113));
 sky130_fd_sc_hd__nand2_2 c141 (.A(net111),
    .B(net943),
    .Y(net114));
 sky130_fd_sc_hd__nor2_8 c142 (.A(net109),
    .B(net113),
    .Y(net115));
 sky130_fd_sc_hd__or2_1 c143 (.A(net114),
    .B(net112),
    .X(net116));
 sky130_fd_sc_hd__nand2_2 c144 (.A(net924),
    .B(net111),
    .Y(net117));
 sky130_fd_sc_hd__and2b_4 c145 (.A_N(net116),
    .B(net1000),
    .X(net118));
 sky130_fd_sc_hd__or3_1 c146 (.A(net115),
    .B(net106),
    .C(net118),
    .X(net119));
 sky130_fd_sc_hd__nor2b_1 c147 (.A(net110),
    .B_N(net118),
    .Y(net120));
 sky130_fd_sc_hd__nand3b_4 c148 (.A_N(net117),
    .B(net107),
    .C(net118),
    .Y(net121));
 sky130_fd_sc_hd__nand3_4 c149 (.A(net113),
    .B(net112),
    .C(net118),
    .Y(net122));
 sky130_fd_sc_hd__or3_4 c150 (.A(net120),
    .B(net921),
    .C(net116),
    .X(net123));
 sky130_fd_sc_hd__or2_4 c151 (.A(net932),
    .B(net122),
    .X(net124));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net120),
    .A1(net124),
    .A2(net122),
    .A3(net108),
    .S0(net107),
    .S1(net935),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 c153 (.A0(net119),
    .A1(net121),
    .A2(net124),
    .A3(net125),
    .S0(net107),
    .S1(net939),
    .X(net126));
 sky130_fd_sc_hd__nand2b_2 c154 (.A_N(net107),
    .B(net928),
    .Y(net127));
 sky130_fd_sc_hd__or2_1 c155 (.A(net15),
    .B(net6),
    .X(net128));
 sky130_fd_sc_hd__nor2_1 c156 (.A(net126),
    .B(net18),
    .Y(net129));
 sky130_fd_sc_hd__nand2_1 c157 (.A(net929),
    .B(net115),
    .Y(net130));
 sky130_fd_sc_hd__and2b_2 c158 (.A_N(net0),
    .B(net115),
    .X(net131));
 sky130_fd_sc_hd__and2_1 c159 (.A(net931),
    .B(net116),
    .X(net132));
 sky130_fd_sc_hd__and2_2 c160 (.A(net928),
    .B(net929),
    .X(net133));
 sky130_fd_sc_hd__or4bb_4 c161 (.A(net132),
    .B(net121),
    .C_N(net0),
    .D_N(net13),
    .X(net134));
 sky130_fd_sc_hd__or2b_4 c162 (.A(net6),
    .B_N(net116),
    .X(net135));
 sky130_fd_sc_hd__nor2b_1 c163 (.A(net988),
    .B_N(net992),
    .Y(net136));
 sky130_fd_sc_hd__or2_4 c164 (.A(net134),
    .B(net13),
    .X(net137));
 sky130_fd_sc_hd__nor2b_1 c165 (.A(net132),
    .B_N(net134),
    .Y(net138));
 sky130_fd_sc_hd__nor2_4 c166 (.A(net128),
    .B(net135),
    .Y(net139));
 sky130_fd_sc_hd__nand2b_1 c167 (.A_N(net129),
    .B(net133),
    .Y(net140));
 sky130_fd_sc_hd__mux4_1 c168 (.A0(net116),
    .A1(net3),
    .A2(net137),
    .A3(net992),
    .S0(net132),
    .S1(net128),
    .X(net141));
 sky130_fd_sc_hd__and2_1 c169 (.A(net140),
    .B(net132),
    .X(net142));
 sky130_fd_sc_hd__or4bb_1 c170 (.A(net110),
    .B(net106),
    .C_N(net142),
    .D_N(net18),
    .X(net143));
 sky130_fd_sc_hd__or4bb_4 c171 (.A(net141),
    .B(net127),
    .C_N(net142),
    .D_N(net107),
    .X(net144));
 sky130_fd_sc_hd__a2111o_1 c172 (.A1(net142),
    .A2(net112),
    .B1(net127),
    .C1(net118),
    .D1(net992),
    .X(net145));
 sky130_fd_sc_hd__a2111oi_4 c173 (.A1(net133),
    .A2(net142),
    .B1(net144),
    .C1(net135),
    .D1(net139),
    .Y(net146));
 sky130_fd_sc_hd__mux4_2 c174 (.A0(net145),
    .A1(net6),
    .A2(net110),
    .A3(net922),
    .S0(net140),
    .S1(net943),
    .X(net147));
 sky130_fd_sc_hd__sdfrbp_2 c175 (.CLK(clknet_4_0_0_clk),
    .D(net138),
    .RESET_B(net144),
    .SCD(net977),
    .SCE(net113),
    .Q(net149),
    .Q_N(net148));
 sky130_fd_sc_hd__or2b_1 c176 (.A(net127),
    .B_N(net25),
    .X(net150));
 sky130_fd_sc_hd__nand2_1 c177 (.A(net27),
    .B(net7),
    .Y(net151));
 sky130_fd_sc_hd__or4bb_1 c178 (.A(net7),
    .B(net25),
    .C_N(net30),
    .D_N(net143),
    .X(net152));
 sky130_fd_sc_hd__and2_1 c179 (.A(net123),
    .B(net134),
    .X(net153));
 sky130_fd_sc_hd__clkinv_16 c187_3 (.A(clknet_1_1__leaf_net898),
    .Y(net1003));
 sky130_fd_sc_hd__or2_1 c181 (.A(net987),
    .B(net23),
    .X(net155));
 sky130_fd_sc_hd__nand2b_1 c182 (.A_N(net21),
    .B(net987),
    .Y(net156));
 sky130_fd_sc_hd__or2_1 c183 (.A(net151),
    .B(net987),
    .X(net157));
 sky130_fd_sc_hd__and2b_1 c184 (.A_N(net3),
    .B(net136),
    .X(net158));
 sky130_fd_sc_hd__sdfbbn_1 c185 (.CLK_N(clknet_4_0_0_clk),
    .D(net36),
    .RESET_B(net143),
    .SCD(net20),
    .SCE(net987),
    .SET_B(net977),
    .Q(net160),
    .Q_N(net159));
 sky130_fd_sc_hd__or2_1 c186 (.A(net158),
    .B(net155),
    .X(net161));
 sky130_fd_sc_hd__inv_1 c344_8 (.A(net918),
    .Y(net1008));
 sky130_fd_sc_hd__and2b_1 c188 (.A_N(net3),
    .B(net160),
    .X(net163));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net161),
    .A1(net156),
    .A2(net158),
    .A3(net139),
    .S0(net3),
    .S1(net153),
    .X(net164));
 sky130_fd_sc_hd__nand2b_1 c190 (.A_N(net150),
    .B(net1002),
    .Y(net165));
 sky130_fd_sc_hd__or4bb_4 c191 (.A(net161),
    .B(net31),
    .C_N(net1007),
    .D_N(net987),
    .X(net166));
 sky130_fd_sc_hd__nor2b_1 c192 (.A(net1001),
    .B_N(net113),
    .Y(net167));
 sky130_fd_sc_hd__a2111oi_0 c193 (.A1(net150),
    .A2(net164),
    .B1(net1006),
    .C1(net9),
    .D1(net987),
    .Y(net168));
 sky130_fd_sc_hd__a2111o_1 c194 (.A1(net160),
    .A2(clknet_1_0__leaf_net168),
    .B1(net161),
    .C1(net30),
    .D1(net974),
    .X(net169));
 sky130_fd_sc_hd__and2b_4 c195 (.A_N(net156),
    .B(clknet_1_0__leaf_net167),
    .X(net170));
 sky130_fd_sc_hd__o2111a_4 c196 (.A1(clknet_1_0__leaf_net165),
    .A2(clknet_1_0__leaf_net170),
    .B1(net107),
    .C1(net158),
    .D1(net776),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net28),
    .A1(net161),
    .A2(net159),
    .A3(net36),
    .S0(clknet_1_0__leaf_net171),
    .X(net172));
 sky130_fd_sc_hd__buf_2 c198 (.A(net731),
    .X(net173));
 sky130_fd_sc_hd__nor2b_2 c199 (.A(net25),
    .B_N(net22),
    .Y(net174));
 sky130_fd_sc_hd__and3b_2 c200 (.A_N(net136),
    .B(net157),
    .C(net174),
    .X(net175));
 sky130_fd_sc_hd__and2b_2 c201 (.A_N(net106),
    .B(net136),
    .X(net176));
 sky130_fd_sc_hd__nor2_1 c202 (.A(net173),
    .B(net49),
    .Y(net177));
 sky130_fd_sc_hd__or4bb_1 c203 (.A(net7),
    .B(net174),
    .C_N(net173),
    .D_N(net148),
    .X(net178));
 sky130_fd_sc_hd__nand3b_4 c204 (.A_N(net157),
    .B(net176),
    .C(net137),
    .Y(net179));
 sky130_fd_sc_hd__buf_1 c205 (.A(net731),
    .X(net180));
 sky130_fd_sc_hd__sdfbbn_1 c206 (.CLK_N(clknet_4_2_0_clk),
    .D(net155),
    .RESET_B(net174),
    .SCD(net1005),
    .SCE(net23),
    .SET_B(net147),
    .Q(net182),
    .Q_N(net181));
 sky130_fd_sc_hd__nand2b_2 c207 (.A_N(net113),
    .B(net157),
    .Y(net183));
 sky130_fd_sc_hd__inv_6 c208 (.A(net915),
    .Y(net184));
 sky130_fd_sc_hd__and2_1 c209 (.A(net182),
    .B(net136),
    .X(net185));
 sky130_fd_sc_hd__mux4_2 c210 (.A0(net23),
    .A1(net182),
    .A2(net184),
    .A3(net185),
    .S0(net136),
    .S1(net987),
    .X(net186));
 sky130_fd_sc_hd__or4bb_2 c211 (.A(net185),
    .B(net186),
    .C_N(net174),
    .D_N(net23),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(net977),
    .A1(net185),
    .A2(net183),
    .A3(net179),
    .S0(net23),
    .S1(net987),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net178),
    .A1(net56),
    .A2(net175),
    .A3(net181),
    .S0(net106),
    .S1(net180),
    .X(net189));
 sky130_fd_sc_hd__nor3b_1 c214 (.A(net135),
    .B(net185),
    .C_N(net820),
    .Y(net190));
 sky130_fd_sc_hd__sdfbbp_1 c215 (.CLK(clknet_4_8_0_clk),
    .D(net180),
    .RESET_B(net190),
    .SCD(net187),
    .SCE(net179),
    .SET_B(net164),
    .Q(net192),
    .Q_N(net191));
 sky130_fd_sc_hd__o2111a_1 c216 (.A1(net59),
    .A2(net180),
    .B1(net186),
    .C1(net181),
    .D1(net820),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net135),
    .A1(net937),
    .A2(net928),
    .A3(net192),
    .S0(net48),
    .S1(net193),
    .X(net194));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net48),
    .A1(net930),
    .A2(net186),
    .A3(net190),
    .S0(net25),
    .S1(net820),
    .X(net195));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net195),
    .A1(net176),
    .A2(net174),
    .A3(net775),
    .S0(net792),
    .S1(net820),
    .X(net196));
 sky130_fd_sc_hd__nand2b_1 c220 (.A_N(net939),
    .B(net19),
    .Y(net197));
 sky130_fd_sc_hd__nand2_2 c221 (.A(net180),
    .B(clknet_1_0__leaf_net170),
    .Y(net198));
 sky130_fd_sc_hd__and3b_1 c222 (.A_N(net57),
    .B(net144),
    .C(net191),
    .X(net199));
 sky130_fd_sc_hd__or2_1 c223 (.A(net186),
    .B(net83),
    .X(net200));
 sky130_fd_sc_hd__nor2_1 c224 (.A(net190),
    .B(net107),
    .Y(net201));
 sky130_fd_sc_hd__nand3_2 c225 (.A(net137),
    .B(net71),
    .C(clknet_1_0__leaf_net198),
    .Y(net202));
 sky130_fd_sc_hd__nand2b_1 c226 (.A_N(net178),
    .B(net78),
    .Y(net203));
 sky130_fd_sc_hd__clkinv_8 c227 (.A(net726),
    .Y(net204));
 sky130_fd_sc_hd__nand2b_2 c228 (.A_N(clknet_1_1__leaf_net170),
    .B(net137),
    .Y(net205));
 sky130_fd_sc_hd__clkbuf_2 c229 (.A(net910),
    .X(net206));
 sky130_fd_sc_hd__or3b_2 c230 (.A(net81),
    .B(net186),
    .C_N(clknet_1_0__leaf_net205),
    .X(net207));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(clknet_1_1__leaf_net202),
    .A1(net204),
    .A2(net985),
    .A3(net191),
    .S0(net83),
    .S1(net206),
    .X(net208));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net206),
    .A1(clknet_1_0__leaf_net208),
    .A2(clknet_1_0__leaf_net207),
    .A3(net204),
    .S0(net985),
    .S1(net144),
    .X(net209));
 sky130_fd_sc_hd__and2_4 c233 (.A(clknet_1_1__leaf_net207),
    .B(net800),
    .X(net210));
 sky130_fd_sc_hd__nand2_4 c234 (.A(clknet_1_1__leaf_net207),
    .B(net985),
    .Y(net211));
 sky130_fd_sc_hd__mux4_2 c235 (.A0(net61),
    .A1(net50),
    .A2(net200),
    .A3(net78),
    .S0(clknet_1_0__leaf_net207),
    .S1(net107),
    .X(net212));
 sky130_fd_sc_hd__nand2b_4 c236 (.A_N(net107),
    .B(clknet_1_0__leaf_net202),
    .Y(net213));
 sky130_fd_sc_hd__clkinv_8 c237 (.A(net726),
    .Y(net214));
 sky130_fd_sc_hd__buf_4 c238 (.A(net910),
    .X(net215));
 sky130_fd_sc_hd__o2111ai_1 c239 (.A1(net49),
    .A2(net206),
    .B1(net214),
    .C1(net187),
    .D1(net82),
    .Y(net216));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net78),
    .A1(net216),
    .A2(net215),
    .A3(net82),
    .S0(net206),
    .S1(net79),
    .X(net217));
 sky130_fd_sc_hd__a2111o_1 c241 (.A1(net199),
    .A2(net206),
    .B1(net215),
    .C1(net214),
    .D1(net985),
    .X(net218));
 sky130_fd_sc_hd__and3_2 c242 (.A(net992),
    .B(net192),
    .C(net787),
    .X(net219));
 sky130_fd_sc_hd__or4bb_4 c243 (.A(net88),
    .B(net85),
    .C_N(net214),
    .D_N(net219),
    .X(net220));
 sky130_fd_sc_hd__or3_2 c244 (.A(net75),
    .B(net941),
    .C(net818),
    .X(net221));
 sky130_fd_sc_hd__and3b_1 c245 (.A_N(net82),
    .B(net814),
    .C(net816),
    .X(net222));
 sky130_fd_sc_hd__nand3_2 c246 (.A(net95),
    .B(net1004),
    .C(net22),
    .Y(net223));
 sky130_fd_sc_hd__inv_1 c247 (.A(net894),
    .Y(net224));
 sky130_fd_sc_hd__or4bb_1 c248 (.A(net52),
    .B(net192),
    .C_N(net22),
    .D_N(net787),
    .X(net225));
 sky130_fd_sc_hd__or3_2 c249 (.A(net222),
    .B(net985),
    .C(net816),
    .X(net226));
 sky130_fd_sc_hd__or2_1 c25 (.A(net923),
    .B(net937),
    .X(net0));
 sky130_fd_sc_hd__or4bb_2 c250 (.A(net92),
    .B(net52),
    .C_N(net992),
    .D_N(net219),
    .X(net227));
 sky130_fd_sc_hd__o2111ai_1 c251 (.A1(net219),
    .A2(net226),
    .B1(net100),
    .C1(net115),
    .D1(net800),
    .Y(net228));
 sky130_fd_sc_hd__sdfrbp_1 c252 (.CLK(clknet_4_10_0_clk),
    .D(net226),
    .RESET_B(net1024),
    .SCD(net1019),
    .SCE(net818),
    .Q(net230),
    .Q_N(net229));
 sky130_fd_sc_hd__sdfbbn_2 c253 (.CLK_N(clknet_4_10_0_clk),
    .D(net224),
    .RESET_B(net82),
    .SCD(net219),
    .SCE(net974),
    .SET_B(net88),
    .Q(net232),
    .Q_N(net231));
 sky130_fd_sc_hd__mux4_4 c254 (.A0(net230),
    .A1(clknet_1_1__leaf_net223),
    .A2(net192),
    .A3(net95),
    .S0(net66),
    .S1(net231),
    .X(net233));
 sky130_fd_sc_hd__or4bb_1 c255 (.A(net52),
    .B(net226),
    .C_N(net232),
    .D_N(net819),
    .X(net234));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net50),
    .A1(net229),
    .A2(net992),
    .A3(net231),
    .S0(net955),
    .S1(net985),
    .X(net235));
 sky130_fd_sc_hd__or4bb_1 c257 (.A(net22),
    .B(net219),
    .C_N(net82),
    .D_N(net203),
    .X(net236));
 sky130_fd_sc_hd__nor3b_1 c258 (.A(net100),
    .B(net235),
    .C_N(net232),
    .Y(net237));
 sky130_fd_sc_hd__a2111oi_2 c259 (.A1(clknet_1_0__leaf_net223),
    .A2(net232),
    .B1(net219),
    .C1(net224),
    .D1(net817),
    .Y(net238));
 sky130_fd_sc_hd__and2_1 c26 (.A(net945),
    .B(net931),
    .X(net1));
 sky130_fd_sc_hd__or4bb_1 c260 (.A(net82),
    .B(net232),
    .C_N(net1019),
    .D_N(net1030),
    .X(net239));
 sky130_fd_sc_hd__or4bb_1 c261 (.A(net219),
    .B(net1000),
    .C_N(net154),
    .D_N(net231),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 c262 (.A(net894),
    .X(net241));
 sky130_fd_sc_hd__sdfbbn_1 c263 (.CLK_N(clknet_4_10_0_clk),
    .D(net101),
    .RESET_B(net226),
    .SCD(net173),
    .SCE(net231),
    .SET_B(net85),
    .Q(net243),
    .Q_N(net242));
 sky130_fd_sc_hd__nor2b_4 c264 (.A(net109),
    .B_N(net117),
    .Y(net244));
 sky130_fd_sc_hd__nor2_1 c265 (.A(net939),
    .B(net934),
    .Y(net245));
 sky130_fd_sc_hd__nand2_4 c266 (.A(net121),
    .B(net939),
    .Y(net948));
 sky130_fd_sc_hd__or2b_2 c267 (.A(net921),
    .B_N(net111),
    .X(net246));
 sky130_fd_sc_hd__or2_2 c268 (.A(net117),
    .B(net245),
    .X(net247));
 sky130_fd_sc_hd__nor2_2 c269 (.A(net119),
    .B(net246),
    .Y(net248));
 sky130_fd_sc_hd__nand2_2 c27 (.A(net940),
    .B(net932),
    .Y(net2));
 sky130_fd_sc_hd__nor2_8 c270 (.A(net124),
    .B(net244),
    .Y(net249));
 sky130_fd_sc_hd__and2_1 c271 (.A(net245),
    .B(net990),
    .X(net250));
 sky130_fd_sc_hd__nand3b_1 c272 (.A_N(net250),
    .B(net989),
    .C(net990),
    .Y(net251));
 sky130_fd_sc_hd__or2b_1 c273 (.A(net990),
    .B_N(net989),
    .X(net252));
 sky130_fd_sc_hd__or3b_4 c274 (.A(net123),
    .B(net942),
    .C_N(net252),
    .X(net253));
 sky130_fd_sc_hd__nand3b_4 c275 (.A_N(net247),
    .B(net253),
    .C(net124),
    .Y(net254));
 sky130_fd_sc_hd__nand2b_1 c276 (.A_N(net246),
    .B(net921),
    .Y(net255));
 sky130_fd_sc_hd__or4bb_4 c277 (.A(net252),
    .B(net245),
    .C_N(net247),
    .D_N(net1000),
    .X(net256));
 sky130_fd_sc_hd__or3b_2 c278 (.A(net111),
    .B(net255),
    .C_N(net256),
    .X(net257));
 sky130_fd_sc_hd__nand2b_2 c279 (.A_N(net255),
    .B(net249),
    .Y(net258));
 sky130_fd_sc_hd__nand2b_2 c28 (.A_N(net945),
    .B(net1),
    .Y(net3));
 sky130_fd_sc_hd__a2111o_2 c280 (.A1(net930),
    .A2(net931),
    .B1(net258),
    .C1(net257),
    .D1(net990),
    .X(net259));
 sky130_fd_sc_hd__mux4_2 c281 (.A0(net245),
    .A1(net257),
    .A2(net250),
    .A3(net252),
    .S0(net124),
    .S1(net246),
    .X(net260));
 sky130_fd_sc_hd__or2_1 c282 (.A(net246),
    .B(net257),
    .X(net261));
 sky130_fd_sc_hd__mux4_2 c283 (.A0(net258),
    .A1(net254),
    .A2(net927),
    .A3(net260),
    .S0(net123),
    .S1(net124),
    .X(net262));
 sky130_fd_sc_hd__mux4_4 c284 (.A0(net255),
    .A1(net259),
    .A2(net244),
    .A3(net262),
    .S0(net111),
    .S1(net124),
    .X(net263));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net263),
    .A1(net260),
    .A2(net1000),
    .A3(net258),
    .S0(net262),
    .S1(net252),
    .X(net264));
 sky130_fd_sc_hd__nor3_1 c286 (.A(net126),
    .B(net139),
    .C(net256),
    .Y(net265));
 sky130_fd_sc_hd__nand2b_1 c287 (.A_N(net258),
    .B(net260),
    .Y(net266));
 sky130_fd_sc_hd__and3b_2 c288 (.A_N(net251),
    .B(net256),
    .C(net989),
    .X(net267));
 sky130_fd_sc_hd__nor2b_2 c289 (.A(net250),
    .B_N(net139),
    .Y(net268));
 sky130_fd_sc_hd__and2_1 c29 (.A(net8),
    .B(net2),
    .X(net4));
 sky130_fd_sc_hd__or3_4 c290 (.A(net265),
    .B(net130),
    .C(net268),
    .X(net269));
 sky130_fd_sc_hd__and2_1 c291 (.A(net927),
    .B(net130),
    .X(net270));
 sky130_fd_sc_hd__or3b_1 c292 (.A(net991),
    .B(net14),
    .C_N(net269),
    .X(net271));
 sky130_fd_sc_hd__o2111a_1 c293 (.A1(net269),
    .A2(net271),
    .B1(net991),
    .C1(net267),
    .D1(net266),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 c294 (.A(net810),
    .X(net273));
 sky130_fd_sc_hd__and2_1 c295 (.A(net244),
    .B(net991),
    .X(net274));
 sky130_fd_sc_hd__nor3_2 c296 (.A(net271),
    .B(net244),
    .C(net269),
    .Y(net275));
 sky130_fd_sc_hd__nand3b_2 c297 (.A_N(net260),
    .B(net130),
    .C(net991),
    .Y(net276));
 sky130_fd_sc_hd__and3b_1 c298 (.A_N(net273),
    .B(net9),
    .C(net276),
    .X(net277));
 sky130_fd_sc_hd__or4bb_1 c299 (.A(net274),
    .B(net13),
    .C_N(net986),
    .D_N(net269),
    .X(net278));
 sky130_fd_sc_hd__or2b_2 c30 (.A(net4),
    .B_N(net1),
    .X(net5));
 sky130_fd_sc_hd__a2111oi_2 c300 (.A1(net278),
    .A2(net269),
    .B1(net139),
    .C1(net276),
    .D1(net991),
    .Y(net279));
 sky130_fd_sc_hd__nor3_2 c301 (.A(net272),
    .B(net275),
    .C(net277),
    .Y(net280));
 sky130_fd_sc_hd__nor3_1 c302 (.A(net121),
    .B(net277),
    .C(net939),
    .Y(net281));
 sky130_fd_sc_hd__mux4_2 c303 (.A0(net267),
    .A1(net268),
    .A2(net276),
    .A3(net250),
    .S0(net279),
    .S1(net258),
    .X(net282));
 sky130_fd_sc_hd__or3_1 c304 (.A(net280),
    .B(net980),
    .C(net276),
    .X(net283));
 sky130_fd_sc_hd__or3b_2 c305 (.A(net277),
    .B(net276),
    .C_N(net258),
    .X(net284));
 sky130_fd_sc_hd__buf_16 c306 (.A(net810),
    .X(net285));
 sky130_fd_sc_hd__nor3_1 c307 (.A(net276),
    .B(net144),
    .C(net285),
    .Y(net286));
 sky130_fd_sc_hd__nand2b_1 c308 (.A_N(net163),
    .B(net123),
    .Y(net287));
 sky130_fd_sc_hd__buf_1 c309 (.A(net784),
    .X(net288));
 sky130_fd_sc_hd__nand2_2 c31 (.A(net2),
    .B(net937),
    .Y(net6));
 sky130_fd_sc_hd__and3b_1 c310 (.A_N(net302),
    .B(net297),
    .C(net306),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(net301),
    .A1(net254),
    .A2(net287),
    .A3(net306),
    .S0(net300),
    .S1(net307),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 c312 (.A(net784),
    .X(net291));
 sky130_fd_sc_hd__inv_2 c313 (.A(net904),
    .Y(net292));
 sky130_fd_sc_hd__clkinv_8 c314 (.A(net746),
    .Y(net293));
 sky130_fd_sc_hd__nor2_1 c315 (.A(net285),
    .B(net13),
    .Y(net294));
 sky130_fd_sc_hd__nor2b_2 c316 (.A(net19),
    .B_N(clknet_1_0__leaf_net165),
    .Y(net295));
 sky130_fd_sc_hd__buf_4 c317 (.A(net746),
    .X(net296));
 sky130_fd_sc_hd__buf_6 c318 (.A(net783),
    .X(net297));
 sky130_fd_sc_hd__and2_1 c319 (.A(net31),
    .B(net297),
    .X(net298));
 sky130_fd_sc_hd__nor2_4 c32 (.A(net933),
    .B(net5),
    .Y(net7));
 sky130_fd_sc_hd__buf_4 c320 (.A(net748),
    .X(net299));
 sky130_fd_sc_hd__or2b_2 c321 (.A(net297),
    .B_N(net285),
    .X(net300));
 sky130_fd_sc_hd__or2_2 c322 (.A(net130),
    .B(net26),
    .X(net301));
 sky130_fd_sc_hd__nand3b_1 c323 (.A_N(net294),
    .B(net301),
    .C(net299),
    .Y(net302));
 sky130_fd_sc_hd__nor2_1 c324 (.A(net139),
    .B(net989),
    .Y(net303));
 sky130_fd_sc_hd__nor2_2 c325 (.A(net280),
    .B(clknet_1_1__leaf_net167),
    .Y(net304));
 sky130_fd_sc_hd__nor2_1 c326 (.A(net944),
    .B(net275),
    .Y(net305));
 sky130_fd_sc_hd__nor2b_4 c327 (.A(net301),
    .B_N(net798),
    .Y(net306));
 sky130_fd_sc_hd__inv_6 c328 (.A(net902),
    .Y(net307));
 sky130_fd_sc_hd__nand3_4 c329 (.A(net267),
    .B(net306),
    .C(net297),
    .Y(net308));
 sky130_fd_sc_hd__and2_1 c33 (.A(net940),
    .B(net925),
    .X(net8));
 sky130_fd_sc_hd__and2_2 c330 (.A(net300),
    .B(net184),
    .X(net309));
 sky130_fd_sc_hd__inv_2 c331 (.A(net915),
    .Y(net310));
 sky130_fd_sc_hd__inv_2 c332 (.A(net766),
    .Y(net311));
 sky130_fd_sc_hd__inv_1 c333 (.A(net797),
    .Y(net312));
 sky130_fd_sc_hd__a2111oi_2 c334 (.A1(net122),
    .A2(net941),
    .B1(net184),
    .C1(net300),
    .D1(clknet_1_0__leaf_net295),
    .Y(net313));
 sky130_fd_sc_hd__mux4_4 c335 (.A0(net982),
    .A1(net122),
    .A2(net990),
    .A3(clknet_1_0__leaf_net295),
    .S0(net930),
    .S1(clknet_1_0__leaf_net313),
    .X(net314));
 sky130_fd_sc_hd__or2b_2 c336 (.A(clknet_1_0__leaf_net313),
    .B_N(net300),
    .X(net315));
 sky130_fd_sc_hd__or3_2 c337 (.A(net293),
    .B(net306),
    .C(net775),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_1 c338 (.A(net797),
    .X(net317));
 sky130_fd_sc_hd__nor2b_1 c339 (.A(net317),
    .B_N(net306),
    .Y(net318));
 sky130_fd_sc_hd__nor2_4 c34 (.A(net923),
    .B(net928),
    .Y(net9));
 sky130_fd_sc_hd__nor3_1 c340 (.A(net987),
    .B(net309),
    .C(net122),
    .Y(net319));
 sky130_fd_sc_hd__inv_2 c341 (.A(net917),
    .Y(net320));
 sky130_fd_sc_hd__inv_2 c342 (.A(net908),
    .Y(net321));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net44),
    .A1(net318),
    .A2(clknet_1_1__leaf_net313),
    .A3(net306),
    .S0(clknet_1_0__leaf_net295),
    .S1(net998),
    .X(net322));
 sky130_fd_sc_hd__clkinv_1 c681_10 (.A(clknet_1_1__leaf_net920),
    .Y(net1010));
 sky130_fd_sc_hd__or4bb_4 c345 (.A(net1009),
    .B(net173),
    .C_N(net998),
    .D_N(net249),
    .X(net324));
 sky130_fd_sc_hd__or2b_1 c346 (.A(net312),
    .B_N(net998),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 c347 (.A(net907),
    .X(net326));
 sky130_fd_sc_hd__or3b_4 c348 (.A(net310),
    .B(net1008),
    .C_N(net300),
    .X(net327));
 sky130_fd_sc_hd__nor3b_2 c349 (.A(net196),
    .B(net326),
    .C_N(net998),
    .Y(net328));
 sky130_fd_sc_hd__o2111ai_4 c35 (.A1(net933),
    .A2(net6),
    .B1(net7),
    .C1(net2),
    .D1(net936),
    .Y(net10));
 sky130_fd_sc_hd__buf_1 c350 (.A(net793),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net982),
    .A1(net325),
    .A2(net328),
    .A3(net998),
    .S0(net310),
    .S1(net989),
    .X(net330));
 sky130_fd_sc_hd__nand3b_1 c352 (.A_N(clknet_1_1__leaf_net205),
    .B(net299),
    .C(net988),
    .Y(net331));
 sky130_fd_sc_hd__and3_1 c353 (.A(net197),
    .B(net299),
    .C(net320),
    .X(net332));
 sky130_fd_sc_hd__or3_1 c354 (.A(net215),
    .B(net83),
    .C(net204),
    .X(net333));
 sky130_fd_sc_hd__nand3b_2 c355 (.A_N(net41),
    .B(net293),
    .C(net988),
    .Y(net334));
 sky130_fd_sc_hd__or4bb_1 c356 (.A(net201),
    .B(clknet_1_0__leaf_net327),
    .C_N(net215),
    .D_N(net30),
    .X(net335));
 sky130_fd_sc_hd__and3_1 c357 (.A(net184),
    .B(net187),
    .C(net988),
    .X(net336));
 sky130_fd_sc_hd__nor3b_1 c358 (.A(net332),
    .B(net214),
    .C_N(net979),
    .Y(net337));
 sky130_fd_sc_hd__buf_1 c359 (.A(net728),
    .X(net338));
 sky130_fd_sc_hd__nand3_2 c36 (.A(net8),
    .B(net10),
    .C(net7),
    .Y(net11));
 sky130_fd_sc_hd__sdfrtn_1 c360 (.CLK_N(clknet_4_9_0_clk),
    .D(net335),
    .RESET_B(net329),
    .SCD(net308),
    .SCE(clknet_1_0__leaf_net198),
    .Q(net339));
 sky130_fd_sc_hd__clkbuf_2 c361 (.A(net727),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net187),
    .A1(net334),
    .A2(net83),
    .A3(net149),
    .S0(clknet_1_0__leaf_net331),
    .S1(net990),
    .X(net341));
 sky130_fd_sc_hd__and3_1 c363 (.A(net83),
    .B(net307),
    .C(net332),
    .X(net342));
 sky130_fd_sc_hd__mux4_2 c364 (.A0(net43),
    .A1(clknet_1_0__leaf_net341),
    .A2(net293),
    .A3(net215),
    .S0(net299),
    .S1(net997),
    .X(net343));
 sky130_fd_sc_hd__inv_1 c365 (.A(net908),
    .Y(net344));
 sky130_fd_sc_hd__sdfrtp_4 c366 (.CLK(clknet_4_9_0_clk),
    .D(net307),
    .RESET_B(net340),
    .SCD(clknet_1_1__leaf_net341),
    .SCE(net215),
    .Q(net345));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net329),
    .A1(clknet_1_1__leaf_net213),
    .A2(net997),
    .A3(net339),
    .S0(net340),
    .S1(clknet_1_1__leaf_net295),
    .X(net346));
 sky130_fd_sc_hd__sdfrtp_1 c368 (.CLK(clknet_4_8_0_clk),
    .D(clknet_1_1__leaf_net341),
    .RESET_B(net338),
    .SCD(net30),
    .SCE(net83),
    .Q(net347));
 sky130_fd_sc_hd__mux4_2 c369 (.A0(net299),
    .A1(net347),
    .A2(clknet_1_1__leaf_net327),
    .A3(clknet_1_0__leaf_net208),
    .S0(net41),
    .S1(net799),
    .X(net348));
 sky130_fd_sc_hd__or3b_2 c37 (.A(net2),
    .B(net926),
    .C_N(net11),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(clknet_1_1__leaf_net331),
    .A1(net347),
    .A2(clknet_1_0__leaf_net208),
    .A3(net299),
    .S0(net799),
    .S1(net822),
    .X(net349));
 sky130_fd_sc_hd__mux4_4 c371 (.A0(net342),
    .A1(net345),
    .A2(net347),
    .A3(net334),
    .S0(net822),
    .S1(clknet_1_0__leaf_net823),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net337),
    .A1(net339),
    .A2(net149),
    .A3(net822),
    .S0(clknet_1_1__leaf_net823),
    .S1(clknet_1_0__leaf_net958),
    .X(net351));
 sky130_fd_sc_hd__mux4_2 c373 (.A0(clknet_1_0__leaf_net331),
    .A1(net197),
    .A2(net922),
    .A3(clknet_1_0__leaf_net341),
    .S0(net347),
    .S1(clknet_1_0__leaf_net823),
    .X(net352));
 sky130_fd_sc_hd__nor3b_2 c374 (.A(net225),
    .B(net94),
    .C_N(clknet_1_0__leaf_net824),
    .Y(net353));
 sky130_fd_sc_hd__or4bb_1 c375 (.A(net173),
    .B(net236),
    .C_N(net231),
    .D_N(net821),
    .X(net354));
 sky130_fd_sc_hd__a2111o_4 c376 (.A1(net334),
    .A2(net338),
    .B1(net985),
    .C1(net992),
    .D1(net797),
    .X(net953));
 sky130_fd_sc_hd__and3b_1 c377 (.A_N(net85),
    .B(net241),
    .C(net344),
    .X(net355));
 sky130_fd_sc_hd__nand3_2 c378 (.A(net985),
    .B(net76),
    .C(net345),
    .Y(net356));
 sky130_fd_sc_hd__nor3_1 c379 (.A(net998),
    .B(net953),
    .C(net985),
    .Y(net357));
 sky130_fd_sc_hd__or2b_4 c38 (.A(net5),
    .B_N(net12),
    .X(net13));
 sky130_fd_sc_hd__or4bb_2 c380 (.A(net353),
    .B(net985),
    .C_N(net76),
    .D_N(net231),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 c381 (.A(net893),
    .X(net359));
 sky130_fd_sc_hd__sdfbbp_1 c382 (.CLK(clknet_4_10_0_clk),
    .D(net236),
    .RESET_B(net235),
    .SCD(net308),
    .SCE(net356),
    .SET_B(net239),
    .Q(net361),
    .Q_N(net360));
 sky130_fd_sc_hd__mux4_2 c383 (.A0(net66),
    .A1(clknet_1_0__leaf_net238),
    .A2(net338),
    .A3(net94),
    .S0(net85),
    .S1(clknet_1_1__leaf_net295),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_2 c384 (.A(net892),
    .X(net362));
 sky130_fd_sc_hd__o2111a_1 c385 (.A1(net356),
    .A2(net998),
    .B1(net974),
    .C1(clknet_1_1__leaf_net358),
    .D1(net85),
    .X(net363));
 sky130_fd_sc_hd__or4bb_2 c386 (.A(net94),
    .B(net173),
    .C_N(clknet_1_1__leaf_net358),
    .D_N(net356),
    .X(net966));
 sky130_fd_sc_hd__mux4_2 c387 (.A0(clknet_1_1__leaf_net238),
    .A1(net125),
    .A2(net85),
    .A3(net94),
    .S0(net988),
    .S1(clknet_1_1__leaf_net958),
    .X(net950));
 sky130_fd_sc_hd__o2111ai_1 c388 (.A1(clknet_1_1__leaf_net358),
    .A2(clknet_1_0__leaf_net970),
    .B1(net125),
    .C1(net356),
    .D1(net799),
    .Y(net364));
 sky130_fd_sc_hd__mux4_4 c389 (.A0(net344),
    .A1(net354),
    .A2(net115),
    .A3(clknet_1_0__leaf_net966),
    .S0(net232),
    .S1(clknet_1_0__leaf_net824),
    .X(net365));
 sky130_fd_sc_hd__nand2b_4 c39 (.A_N(net1),
    .B(net10),
    .Y(net14));
 sky130_fd_sc_hd__mux4_4 c390 (.A0(net357),
    .A1(net232),
    .A2(clknet_1_0__leaf_net358),
    .A3(clknet_1_0__leaf_net966),
    .S0(clknet_1_0__leaf_net806),
    .S1(net821),
    .X(net366));
 sky130_fd_sc_hd__mux4_2 c391 (.A0(net239),
    .A1(clknet_1_1__leaf_net233),
    .A2(net66),
    .A3(net953),
    .S0(net989),
    .S1(net828),
    .X(net367));
 sky130_fd_sc_hd__mux4_4 c392 (.A0(net214),
    .A1(net366),
    .A2(clknet_1_0__leaf_net358),
    .A3(net998),
    .S0(net227),
    .S1(net827),
    .X(net368));
 sky130_fd_sc_hd__or4bb_1 c393 (.A(net1000),
    .B(clknet_1_0__leaf_net966),
    .C_N(clknet_1_1__leaf_net824),
    .D_N(net828),
    .X(net369));
 sky130_fd_sc_hd__mux4_2 c394 (.A0(net367),
    .A1(clknet_1_0__leaf_net966),
    .A2(clknet_1_0__leaf_net369),
    .A3(net953),
    .S0(net345),
    .S1(net797),
    .X(net370));
 sky130_fd_sc_hd__sdfrtp_1 c395 (.CLK(clknet_4_11_0_clk),
    .D(net354),
    .RESET_B(clknet_1_1__leaf_net369),
    .SCD(net1027),
    .SCE(net830),
    .Q(net962));
 sky130_fd_sc_hd__nand2_2 c396 (.A(net935),
    .B(net261),
    .Y(net371));
 sky130_fd_sc_hd__nor2b_1 c397 (.A(net125),
    .B_N(net990),
    .Y(net372));
 sky130_fd_sc_hd__and2b_1 c398 (.A_N(net934),
    .B(net935),
    .X(net373));
 sky130_fd_sc_hd__and2_1 c399 (.A(net259),
    .B(net257),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c40 (.A0(net10),
    .A1(net4),
    .A2(net6),
    .A3(net14),
    .S0(net7),
    .S1(net8),
    .X(net15));
 sky130_fd_sc_hd__nor2b_1 c400 (.A(net374),
    .B_N(net941),
    .Y(net375));
 sky130_fd_sc_hd__and2b_1 c401 (.A_N(net373),
    .B(net262),
    .X(net376));
 sky130_fd_sc_hd__nor2_1 c402 (.A(net264),
    .B(net983),
    .Y(net377));
 sky130_fd_sc_hd__and2_1 c403 (.A(net252),
    .B(net375),
    .X(net378));
 sky130_fd_sc_hd__nand2b_4 c404 (.A_N(net378),
    .B(net373),
    .Y(net379));
 sky130_fd_sc_hd__nand2b_1 c405 (.A_N(net257),
    .B(net983),
    .Y(net380));
 sky130_fd_sc_hd__and2_1 c406 (.A(net261),
    .B(net378),
    .X(net381));
 sky130_fd_sc_hd__nand2b_1 c407 (.A_N(net375),
    .B(net262),
    .Y(net382));
 sky130_fd_sc_hd__nand2_1 c408 (.A(net262),
    .B(net380),
    .Y(net383));
 sky130_fd_sc_hd__inv_4 c409 (.A(net811),
    .Y(net384));
 sky130_fd_sc_hd__nand2_2 c41 (.A(net15),
    .B(net936),
    .Y(net16));
 sky130_fd_sc_hd__mux4_1 c410 (.A0(net377),
    .A1(net115),
    .A2(net114),
    .A3(net257),
    .S0(net379),
    .S1(net261),
    .X(net385));
 sky130_fd_sc_hd__buf_6 c411 (.A(net811),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_4 c412 (.A(net899),
    .X(net387));
 sky130_fd_sc_hd__nor2b_4 c413 (.A(net387),
    .B_N(net807),
    .Y(net388));
 sky130_fd_sc_hd__or2b_2 c414 (.A(clknet_1_0__leaf_net388),
    .B_N(net376),
    .X(net389));
 sky130_fd_sc_hd__nor2b_1 c415 (.A(net382),
    .B_N(clknet_1_0__leaf_net389),
    .Y(net390));
 sky130_fd_sc_hd__a2111o_1 c416 (.A1(net374),
    .A2(clknet_1_0__leaf_net390),
    .B1(net381),
    .C1(net983),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_4 c417 (.A(net783),
    .X(net949));
 sky130_fd_sc_hd__nor3b_4 c418 (.A(net943),
    .B(net991),
    .C_N(net268),
    .Y(net392));
 sky130_fd_sc_hd__nand3b_1 c419 (.A_N(net980),
    .B(net983),
    .C(net13),
    .Y(net393));
 sky130_fd_sc_hd__mux4_2 c42 (.A0(net0),
    .A1(net938),
    .A2(net2),
    .A3(net988),
    .S0(net13),
    .S1(net12),
    .X(net17));
 sky130_fd_sc_hd__nor3b_2 c420 (.A(net149),
    .B(net980),
    .C_N(net983),
    .Y(net394));
 sky130_fd_sc_hd__buf_2 c421 (.A(clknet_1_0__leaf_net897),
    .X(net395));
 sky130_fd_sc_hd__nand3_1 c422 (.A(net937),
    .B(net256),
    .C(net983),
    .Y(net396));
 sky130_fd_sc_hd__a2111o_1 c423 (.A1(net378),
    .A2(net384),
    .B1(net268),
    .C1(net1000),
    .D1(net990),
    .X(net397));
 sky130_fd_sc_hd__dlymetal6s2s_1 c424 (.A(clknet_1_1__leaf_net897),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_2 c425 (.A(net905),
    .X(net399));
 sky130_fd_sc_hd__sdfbbn_1 c426 (.CLK_N(clknet_4_1_0_clk),
    .D(net384),
    .RESET_B(net379),
    .SCD(net135),
    .SCE(net392),
    .SET_B(clknet_1_0__leaf_net395),
    .Q(net401),
    .Q_N(net400));
 sky130_fd_sc_hd__and3b_1 c427 (.A_N(net375),
    .B(net396),
    .C(net269),
    .X(net402));
 sky130_fd_sc_hd__and3b_4 c428 (.A_N(net392),
    .B(net402),
    .C(net400),
    .X(net959));
 sky130_fd_sc_hd__sdfsbp_1 c429 (.CLK(clknet_4_1_0_clk),
    .D(net941),
    .SCD(net959),
    .SCE(net983),
    .SET_B(net1021),
    .Q(net404),
    .Q_N(net403));
 sky130_fd_sc_hd__or4bb_2 c43 (.A(net13),
    .B(net12),
    .C_N(net17),
    .D_N(net15),
    .X(net18));
 sky130_fd_sc_hd__mux4_4 c430 (.A0(net402),
    .A1(clknet_1_0__leaf_net398),
    .A2(net399),
    .A3(net403),
    .S0(net266),
    .S1(net375),
    .X(net405));
 sky130_fd_sc_hd__o2111a_4 c431 (.A1(clknet_1_0__leaf_net395),
    .A2(net392),
    .B1(net403),
    .C1(net379),
    .D1(net118),
    .X(net406));
 sky130_fd_sc_hd__o2111a_4 c432 (.A1(clknet_1_0__leaf_net405),
    .A2(net247),
    .B1(net399),
    .C1(net992),
    .D1(clknet_1_0__leaf_net390),
    .X(net407));
 sky130_fd_sc_hd__mux4_2 c433 (.A0(net266),
    .A1(net127),
    .A2(net983),
    .A3(net959),
    .S0(clknet_1_0__leaf_net398),
    .S1(net804),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net376),
    .A1(net991),
    .A2(net393),
    .A3(net959),
    .S0(net269),
    .S1(net831),
    .X(net409));
 sky130_fd_sc_hd__mux4_4 c435 (.A0(clknet_1_0__leaf_net405),
    .A1(net935),
    .A2(net393),
    .A3(net269),
    .S0(net979),
    .S1(net832),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net269),
    .A1(clknet_1_1__leaf_net398),
    .A2(clknet_1_1__leaf_net405),
    .A3(net270),
    .S0(net147),
    .S1(net833),
    .X(net411));
 sky130_fd_sc_hd__or3_2 c437 (.A(net404),
    .B(net815),
    .C(net833),
    .X(net412));
 sky130_fd_sc_hd__nor3_2 c438 (.A(net399),
    .B(net404),
    .C(net833),
    .Y(net413));
 sky130_fd_sc_hd__mux4_4 c439 (.A0(net396),
    .A1(clknet_1_1__leaf_net405),
    .A2(clknet_1_0__leaf_net390),
    .A3(net996),
    .S1(net832),
    .X(net414));
 sky130_fd_sc_hd__and2_4 c44 (.A(net5),
    .B(net40),
    .X(net19));
 sky130_fd_sc_hd__nor2_4 c440 (.A(clknet_1_1__leaf_net395),
    .B(net803),
    .Y(net415));
 sky130_fd_sc_hd__nor2b_4 c441 (.A(net415),
    .B_N(net936),
    .Y(net416));
 sky130_fd_sc_hd__nor2b_1 c442 (.A(net287),
    .B_N(net117),
    .Y(net417));
 sky130_fd_sc_hd__or3b_4 c443 (.A(net268),
    .B(clknet_1_1__leaf_net167),
    .C_N(net20),
    .X(net418));
 sky130_fd_sc_hd__or3b_4 c444 (.A(clknet_1_0__leaf_net416),
    .B(net9),
    .C_N(net979),
    .X(net419));
 sky130_fd_sc_hd__or2b_4 c445 (.A(net296),
    .B_N(net832),
    .X(net420));
 sky130_fd_sc_hd__nor3b_1 c446 (.A(net20),
    .B(net135),
    .C_N(net420),
    .Y(net421));
 sky130_fd_sc_hd__nand2_4 c447 (.A(net288),
    .B(clknet_1_1__leaf_net165),
    .Y(net422));
 sky130_fd_sc_hd__clkbuf_1 c448 (.A(net747),
    .X(net423));
 sky130_fd_sc_hd__a2111o_1 c449 (.A1(net305),
    .A2(net268),
    .B1(clknet_1_0__leaf_net390),
    .C1(clknet_1_0__leaf_net422),
    .D1(net386),
    .X(net424));
 sky130_fd_sc_hd__and2_2 c45 (.A(net925),
    .B(net40),
    .X(net20));
 sky130_fd_sc_hd__or4bb_1 c450 (.A(net423),
    .B(net19),
    .C_N(clknet_1_0__leaf_net416),
    .D_N(net420),
    .X(net425));
 sky130_fd_sc_hd__o2111ai_1 c451 (.A1(clknet_1_1__leaf_net422),
    .A2(net983),
    .B1(net403),
    .C1(net256),
    .D1(net815),
    .Y(net426));
 sky130_fd_sc_hd__or4bb_1 c452 (.A(clknet_1_0__leaf_net425),
    .B(net292),
    .C_N(net256),
    .D_N(net832),
    .X(net427));
 sky130_fd_sc_hd__and2_1 c453 (.A(net417),
    .B(clknet_1_0__leaf_net426),
    .X(net428));
 sky130_fd_sc_hd__or2b_1 c454 (.A(net427),
    .B_N(net420),
    .X(net429));
 sky130_fd_sc_hd__nor2_4 c455 (.A(clknet_1_0__leaf_net428),
    .B(net420),
    .Y(net430));
 sky130_fd_sc_hd__nor3b_4 c456 (.A(net404),
    .B(clknet_1_1__leaf_net416),
    .C_N(net420),
    .Y(net431));
 sky130_fd_sc_hd__and2_2 c457 (.A(net429),
    .B(net831),
    .X(net432));
 sky130_fd_sc_hd__nor2_1 c458 (.A(net936),
    .B(net786),
    .Y(net433));
 sky130_fd_sc_hd__mux4_4 c459 (.A0(net144),
    .A1(clknet_1_1__leaf_net430),
    .A2(clknet_1_0__leaf_net428),
    .A3(net433),
    .S0(net20),
    .S1(net941),
    .X(net434));
 sky130_fd_sc_hd__nand2b_1 c46 (.A_N(net927),
    .B(net925),
    .Y(net21));
 sky130_fd_sc_hd__mux4_4 c460 (.A0(net418),
    .A1(net413),
    .A2(net986),
    .A3(clknet_1_1__leaf_net425),
    .S0(net988),
    .S1(net999),
    .X(net435));
 sky130_fd_sc_hd__mux4_4 c461 (.A0(net433),
    .A1(net959),
    .A2(clknet_1_1__leaf_net428),
    .A3(clknet_1_0__leaf_net435),
    .S0(net420),
    .S1(net999),
    .X(net436));
 sky130_fd_sc_hd__or4bb_4 c462 (.A(clknet_1_1__leaf_net390),
    .B(net309),
    .C_N(net328),
    .D_N(net183),
    .X(net437));
 sky130_fd_sc_hd__buf_16 c463 (.A(net895),
    .X(net438));
 sky130_fd_sc_hd__buf_16 c464 (.A(net895),
    .X(net439));
 sky130_fd_sc_hd__inv_4 c465 (.A(net901),
    .Y(net440));
 sky130_fd_sc_hd__mux4_4 c466 (.A0(net183),
    .A1(net401),
    .A2(net997),
    .A3(clknet_1_1__leaf_net390),
    .S0(net942),
    .S1(net249),
    .X(net441));
 sky130_fd_sc_hd__nand3b_4 c467 (.A_N(net438),
    .B(net946),
    .C(net792),
    .Y(net442));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(clknet_1_0__leaf_net171),
    .A1(clknet_1_0__leaf_net432),
    .A2(net996),
    .A3(net293),
    .S1(net791),
    .X(net443));
 sky130_fd_sc_hd__buf_16 c469 (.A(net900),
    .X(net444));
 sky130_fd_sc_hd__and2b_4 c47 (.A_N(net925),
    .B(net938),
    .X(net22));
 sky130_fd_sc_hd__sdfsbp_1 c470 (.CLK(clknet_4_3_0_clk),
    .D(net179),
    .SCD(net293),
    .SCE(net815),
    .SET_B(net999),
    .Q(net445));
 sky130_fd_sc_hd__nor3b_4 c471 (.A(clknet_1_1__leaf_net398),
    .B(net442),
    .C_N(net936),
    .Y(net446));
 sky130_fd_sc_hd__nor3b_1 c472 (.A(net249),
    .B(net979),
    .C_N(net781),
    .Y(net447));
 sky130_fd_sc_hd__sdfstp_1 c473 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net165),
    .SCD(clknet_1_0__leaf_net432),
    .SCE(net447),
    .SET_B(net444),
    .Q(net448));
 sky130_fd_sc_hd__clkinv_4 c474 (.A(net767),
    .Y(net449));
 sky130_fd_sc_hd__nor3_2 c475 (.A(net306),
    .B(net989),
    .C(net941),
    .Y(net450));
 sky130_fd_sc_hd__sdfbbn_2 c476 (.CLK_N(clknet_4_12_0_clk),
    .D(net309),
    .RESET_B(net976),
    .SCD(net448),
    .SCE(clknet_1_0__leaf_net446),
    .SET_B(net983),
    .Q(net452),
    .Q_N(net451));
 sky130_fd_sc_hd__mux4_2 c477 (.A0(net442),
    .A1(net328),
    .A2(net448),
    .A3(net976),
    .S0(clknet_1_0__leaf_net430),
    .S1(net386),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net438),
    .A1(net442),
    .A2(net976),
    .A3(net448),
    .S0(net449),
    .S1(net451),
    .X(net454));
 sky130_fd_sc_hd__mux4_2 c479 (.A0(net992),
    .A1(clknet_1_1__leaf_net430),
    .A2(net449),
    .A3(net448),
    .S0(net999),
    .S1(net838),
    .X(net455));
 sky130_fd_sc_hd__or2_2 c48 (.A(net21),
    .B(net40),
    .X(net23));
 sky130_fd_sc_hd__mux4_4 c480 (.A0(net445),
    .A1(net452),
    .A2(net976),
    .A3(net448),
    .S0(net979),
    .S1(net839),
    .X(net456));
 sky130_fd_sc_hd__mux4_2 c481 (.A0(net448),
    .A1(clknet_1_1__leaf_net432),
    .A2(net254),
    .A3(net831),
    .S0(net839),
    .S1(net840),
    .X(net457));
 sky130_fd_sc_hd__sdfbbp_1 c482 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net432),
    .RESET_B(net452),
    .SCD(net449),
    .SCE(net438),
    .SET_B(net812),
    .Q(net458));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net421),
    .A1(net447),
    .A2(net309),
    .A3(clknet_1_0__leaf_net446),
    .S0(net837),
    .S1(net841),
    .X(net459));
 sky130_fd_sc_hd__sdfbbn_2 c484 (.CLK_N(clknet_4_12_0_clk),
    .D(net394),
    .RESET_B(clknet_1_0__leaf_net198),
    .SCD(net785),
    .SCE(clknet_1_0__leaf_net823),
    .SET_B(net635),
    .Q(net461),
    .Q_N(net460));
 sky130_fd_sc_hd__o2111a_1 c485 (.A1(net293),
    .A2(net979),
    .B1(net248),
    .C1(net936),
    .D1(net825),
    .X(net462));
 sky130_fd_sc_hd__mux4_2 c486 (.A0(net71),
    .A1(net943),
    .A2(net460),
    .A3(net988),
    .S0(clknet_1_0__leaf_net823),
    .S1(net999),
    .X(net463));
 sky130_fd_sc_hd__mux4_4 c487 (.A0(clknet_1_0__leaf_net211),
    .A1(clknet_1_0__leaf_net324),
    .A2(net54),
    .A3(net450),
    .S0(net79),
    .S1(net825),
    .X(net464));
 sky130_fd_sc_hd__sdfbbn_1 c488 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net208),
    .RESET_B(net117),
    .SCD(net293),
    .SCE(net922),
    .SET_B(clknet_1_0__leaf_net958),
    .Q(net466),
    .Q_N(net465));
 sky130_fd_sc_hd__mux4_2 c489 (.A0(net179),
    .A1(net76),
    .A2(net440),
    .A3(clknet_1_0__leaf_net198),
    .S0(net786),
    .S1(net841),
    .X(net467));
 sky130_fd_sc_hd__or2b_1 c49 (.A(net12),
    .B_N(net40),
    .X(net24));
 sky130_fd_sc_hd__sdfbbp_1 c490 (.CLK(clknet_4_14_0_clk),
    .D(net462),
    .RESET_B(net76),
    .SCD(net465),
    .SCE(net450),
    .SET_B(clknet_1_0__leaf_net843),
    .Q(net469),
    .Q_N(net468));
 sky130_fd_sc_hd__a2111o_1 c491 (.A1(net340),
    .A2(net466),
    .B1(net76),
    .C1(net468),
    .D1(net831),
    .X(net470));
 sky130_fd_sc_hd__mux4_4 c492 (.A0(net450),
    .A1(net179),
    .A2(clknet_1_1__leaf_net211),
    .A3(net470),
    .S0(clknet_1_1__leaf_net208),
    .S1(net340),
    .X(net471));
 sky130_fd_sc_hd__o2111ai_2 c493 (.A1(net79),
    .A2(net460),
    .B1(net997),
    .C1(clknet_1_1__leaf_net843),
    .D1(clknet_1_0__leaf_net844),
    .Y(net472));
 sky130_fd_sc_hd__sdfbbn_2 c494 (.CLK_N(clknet_4_12_0_clk),
    .D(net371),
    .RESET_B(net118),
    .SCD(net462),
    .SCE(net959),
    .SET_B(clknet_1_0__leaf_net844),
    .Q(net474),
    .Q_N(net473));
 sky130_fd_sc_hd__a2111oi_0 c495 (.A1(clknet_1_1__leaf_net324),
    .A2(net470),
    .B1(net345),
    .C1(net465),
    .D1(clknet_1_0__leaf_net844),
    .Y(net475));
 sky130_fd_sc_hd__mux4_2 c496 (.A0(net470),
    .A1(clknet_1_0__leaf_net472),
    .A2(net466),
    .A3(net144),
    .S0(net785),
    .S1(clknet_1_0__leaf_net844),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net19),
    .A1(net71),
    .A2(clknet_1_1__leaf_net208),
    .A3(net461),
    .S0(net473),
    .S1(net635),
    .X(net477));
 sky130_fd_sc_hd__a2111oi_1 c498 (.A1(net440),
    .A2(net936),
    .B1(clknet_1_0__leaf_net472),
    .C1(net943),
    .D1(clknet_1_1__leaf_net463),
    .Y(net478));
 sky130_fd_sc_hd__sdfbbn_1 c499 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net476),
    .RESET_B(clknet_1_0__leaf_net478),
    .SCD(net974),
    .SCE(net780),
    .SET_B(net821),
    .Q(net480),
    .Q_N(net479));
 sky130_fd_sc_hd__and2b_2 c50 (.A_N(net9),
    .B(net22),
    .X(net25));
 sky130_fd_sc_hd__sdfbbp_1 c500 (.CLK(clknet_4_14_0_clk),
    .D(net394),
    .RESET_B(net449),
    .SCD(net54),
    .SCE(net470),
    .SET_B(clknet_1_1__leaf_net844),
    .Q(net482),
    .Q_N(net481));
 sky130_fd_sc_hd__mux4_4 c501 (.A0(clknet_1_0__leaf_net478),
    .A1(net481),
    .A2(clknet_1_0__leaf_net476),
    .A3(net974),
    .S0(net460),
    .S1(net780),
    .X(net483));
 sky130_fd_sc_hd__mux4_2 c502 (.A0(net469),
    .A1(clknet_1_0__leaf_net475),
    .A2(net479),
    .A3(net282),
    .S0(net162),
    .S1(net845),
    .X(net484));
 sky130_fd_sc_hd__mux4_4 c503 (.A0(net480),
    .A1(net484),
    .A2(clknet_1_1__leaf_net463),
    .A3(clknet_1_0__leaf_net475),
    .S0(net949),
    .S1(net846),
    .X(net485));
 sky130_fd_sc_hd__mux4_4 c504 (.A0(net482),
    .A1(clknet_1_1__leaf_net475),
    .A2(clknet_1_1__leaf_net478),
    .A3(net821),
    .S0(net845),
    .S1(net848),
    .X(net486));
 sky130_fd_sc_hd__mux4_2 c505 (.A0(net486),
    .A1(clknet_1_1__leaf_net475),
    .A2(clknet_1_1__leaf_net198),
    .A3(clknet_1_1__leaf_net478),
    .S0(net846),
    .S1(net847),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c509 (.A0(net308),
    .A1(clknet_1_1__leaf_net369),
    .A2(net992),
    .A3(clknet_1_1__leaf_net472),
    .S0(net240),
    .S1(clknet_1_0__leaf_net950),
    .X(net488));
 sky130_fd_sc_hd__and2_2 c51 (.A(net24),
    .B(net7),
    .X(net26));
 sky130_fd_sc_hd__mux4_2 c510 (.A0(clknet_1_0__leaf_net472),
    .A1(net953),
    .A2(net221),
    .A3(net955),
    .S0(net231),
    .S1(net131),
    .X(net489));
 sky130_fd_sc_hd__mux4_2 c511 (.A0(net232),
    .A1(net955),
    .A2(clknet_1_1__leaf_net472),
    .A3(clknet_1_0__leaf_net966),
    .S0(clknet_1_0__leaf_net369),
    .S1(clknet_1_1__leaf_net806),
    .X(net490));
 sky130_fd_sc_hd__o2111ai_2 c512 (.A1(net221),
    .A2(net943),
    .B1(net362),
    .C1(net988),
    .D1(clknet_1_1__leaf_net958),
    .Y(net967));
 sky130_fd_sc_hd__mux4_2 c513 (.A0(net243),
    .A1(net240),
    .A2(net939),
    .A3(net220),
    .S0(clknet_1_1__leaf_net472),
    .S1(clknet_1_1__leaf_net966),
    .X(net491));
 sky130_fd_sc_hd__mux4_4 c514 (.A0(net125),
    .A1(net946),
    .A2(net974),
    .A3(net220),
    .S0(clknet_1_1__leaf_net823),
    .S1(clknet_1_1__leaf_net958),
    .X(net492));
 sky130_fd_sc_hd__o2111ai_1 c515 (.A1(net76),
    .A2(net232),
    .B1(net955),
    .C1(net830),
    .D1(net853),
    .Y(net493));
 sky130_fd_sc_hd__sdfbbn_1 c516 (.CLK_N(clknet_4_11_0_clk),
    .D(net227),
    .RESET_B(net220),
    .SCD(net359),
    .SCE(net821),
    .SET_B(net1022),
    .Q(net494));
 sky130_fd_sc_hd__mux4_1 c517 (.A0(net220),
    .A1(clknet_1_1__leaf_net472),
    .A2(clknet_1_1__leaf_net369),
    .A3(clknet_1_1__leaf_net295),
    .S0(net821),
    .S1(net852),
    .X(net495));
 sky130_fd_sc_hd__sdfbbn_1 c518 (.CLK_N(clknet_4_10_0_clk),
    .D(net359),
    .RESET_B(net361),
    .SCD(net1026),
    .SCE(net974),
    .SET_B(clknet_1_1__leaf_net823),
    .Q(net961));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net439),
    .A1(net362),
    .A2(net149),
    .A3(clknet_1_0__leaf_net472),
    .S0(net959),
    .S1(net853),
    .X(net496));
 sky130_fd_sc_hd__or2b_2 c52 (.A(net40),
    .B_N(net20),
    .X(net27));
 sky130_fd_sc_hd__o2111ai_2 c520 (.A1(net345),
    .A2(net162),
    .B1(net955),
    .C1(clknet_1_0__leaf_net369),
    .D1(net959),
    .Y(net497));
 sky130_fd_sc_hd__sdfbbp_1 c521 (.CLK(clknet_4_11_0_clk),
    .D(net131),
    .RESET_B(net355),
    .SCD(net955),
    .SCE(net148),
    .SET_B(clknet_1_1__leaf_net823),
    .Q(net499),
    .Q_N(net498));
 sky130_fd_sc_hd__o2111ai_4 c522 (.A1(net955),
    .A2(net498),
    .B1(net953),
    .C1(net851),
    .D1(net854),
    .Y(net500));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(clknet_1_1__leaf_net295),
    .A1(net974),
    .A2(net500),
    .A3(net498),
    .S0(net959),
    .S1(net162),
    .X(net501));
 sky130_fd_sc_hd__a2111o_4 c524 (.A1(net500),
    .A2(net499),
    .B1(net360),
    .C1(net105),
    .D1(clknet_1_1__leaf_net472),
    .X(net956));
 sky130_fd_sc_hd__mux4_2 c525 (.A0(net499),
    .A1(clknet_1_0__leaf_net956),
    .A2(net500),
    .A3(net989),
    .S0(net812),
    .S1(net853),
    .X(net963));
 sky130_fd_sc_hd__mux4_2 c526 (.A0(net489),
    .A1(net493),
    .A2(clknet_1_1__leaf_net956),
    .A3(clknet_1_1__leaf_net369),
    .S0(net500),
    .S1(net855),
    .X(net502));
 sky130_fd_sc_hd__mux4_4 c527 (.A0(net989),
    .A1(net494),
    .A2(clknet_1_0__leaf_net956),
    .A3(net355),
    .S0(net830),
    .S1(net856),
    .X(net503));
 sky130_fd_sc_hd__nand3_1 c528 (.A(net931),
    .B(net259),
    .C(net944),
    .Y(net504));
 sky130_fd_sc_hd__and2_1 c529 (.A(clknet_1_1__leaf_net388),
    .B(net259),
    .X(net505));
 sky130_fd_sc_hd__nand2_1 c53 (.A(net22),
    .B(net24),
    .Y(net28));
 sky130_fd_sc_hd__buf_2 c530 (.A(net788),
    .X(net506));
 sky130_fd_sc_hd__or2b_1 c531 (.A(net504),
    .B_N(net922),
    .X(net507));
 sky130_fd_sc_hd__or2_2 c532 (.A(net505),
    .B(net114),
    .X(net508));
 sky130_fd_sc_hd__or2b_2 c533 (.A(net372),
    .B_N(net506),
    .X(net509));
 sky130_fd_sc_hd__nor2b_1 c534 (.A(net921),
    .B_N(net256),
    .Y(net510));
 sky130_fd_sc_hd__or2_2 c535 (.A(net510),
    .B(net259),
    .X(net511));
 sky130_fd_sc_hd__and2b_1 c536 (.A_N(net942),
    .B(net509),
    .X(net512));
 sky130_fd_sc_hd__or2_2 c537 (.A(clknet_1_1__leaf_net508),
    .B(net512),
    .X(net513));
 sky130_fd_sc_hd__nor3b_4 c538 (.A(net509),
    .B(net506),
    .C_N(net510),
    .Y(net514));
 sky130_fd_sc_hd__and3_1 c539 (.A(net506),
    .B(net509),
    .C(net934),
    .X(net515));
 sky130_fd_sc_hd__or4bb_1 c54 (.A(net20),
    .B(net27),
    .C_N(net22),
    .D_N(net942),
    .X(net29));
 sky130_fd_sc_hd__a2111oi_2 c540 (.A1(net506),
    .A2(net504),
    .B1(clknet_1_0__leaf_net513),
    .C1(net984),
    .D1(net249),
    .Y(net516));
 sky130_fd_sc_hd__or2_1 c541 (.A(net509),
    .B(net510),
    .X(net517));
 sky130_fd_sc_hd__nand3b_4 c542 (.A_N(net510),
    .B(net372),
    .C(net984),
    .Y(net518));
 sky130_fd_sc_hd__mux4_2 c543 (.A0(net517),
    .A1(net518),
    .A2(net509),
    .A3(clknet_1_0__leaf_net513),
    .S0(net506),
    .S1(clknet_1_0__leaf_net508),
    .X(net519));
 sky130_fd_sc_hd__or3b_1 c544 (.A(net515),
    .B(net944),
    .C_N(net518),
    .X(net520));
 sky130_fd_sc_hd__nand2b_2 c545 (.A_N(net512),
    .B(net511),
    .Y(net521));
 sky130_fd_sc_hd__and3_1 c546 (.A(net380),
    .B(net984),
    .C(net521),
    .X(net522));
 sky130_fd_sc_hd__buf_1 c547 (.A(net788),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net507),
    .A1(net522),
    .A2(clknet_1_0__leaf_net519),
    .A3(net523),
    .S0(net506),
    .S1(net512),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net253),
    .A1(net506),
    .A2(net379),
    .A3(net518),
    .S0(net807),
    .S1(net857),
    .X(net525));
 sky130_fd_sc_hd__and2b_4 c55 (.A_N(net29),
    .B(net21),
    .X(net30));
 sky130_fd_sc_hd__or2b_1 c550 (.A(net991),
    .B_N(net996),
    .X(net526));
 sky130_fd_sc_hd__inv_2 c551 (.A(net779),
    .Y(net527));
 sky130_fd_sc_hd__and2_1 c552 (.A(net284),
    .B(net518),
    .X(net528));
 sky130_fd_sc_hd__or2b_1 c553 (.A(net520),
    .B_N(clknet_1_0__leaf_net513),
    .X(net529));
 sky130_fd_sc_hd__inv_4 c554 (.A(net779),
    .Y(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 c555 (.A(net899),
    .X(net531));
 sky130_fd_sc_hd__nor2b_1 c556 (.A(net18),
    .B_N(net530),
    .Y(net532));
 sky130_fd_sc_hd__inv_2 c557 (.A(net750),
    .Y(net533));
 sky130_fd_sc_hd__nand2b_1 c558 (.A_N(net527),
    .B(net518),
    .Y(net534));
 sky130_fd_sc_hd__and3b_4 c559 (.A_N(net383),
    .B(net523),
    .C(net984),
    .X(net535));
 sky130_fd_sc_hd__and2_1 c56 (.A(net29),
    .B(net28),
    .X(net31));
 sky130_fd_sc_hd__inv_2 c560 (.A(net907),
    .Y(net965));
 sky130_fd_sc_hd__buf_1 c561 (.A(net749),
    .X(net536));
 sky130_fd_sc_hd__buf_1 c562 (.A(net909),
    .X(net537));
 sky130_fd_sc_hd__buf_6 c563 (.A(net906),
    .X(net538));
 sky130_fd_sc_hd__a2111oi_1 c564 (.A1(net134),
    .A2(net532),
    .B1(net284),
    .C1(net115),
    .D1(net521),
    .Y(net539));
 sky130_fd_sc_hd__or4bb_1 c565 (.A(net536),
    .B(clknet_1_0__leaf_net531),
    .C_N(net535),
    .D_N(net990),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net530),
    .A1(net528),
    .A2(net1032),
    .A3(net284),
    .S0(net535),
    .S1(net779),
    .X(net541));
 sky130_fd_sc_hd__mux4_4 c567 (.A0(net538),
    .A1(net536),
    .A2(net535),
    .A3(net530),
    .S0(net991),
    .S1(net949),
    .X(net542));
 sky130_fd_sc_hd__inv_4 c568 (.A(net917),
    .Y(net543));
 sky130_fd_sc_hd__buf_8 c569 (.A(clknet_1_1__leaf_net919),
    .X(net544));
 sky130_fd_sc_hd__or4bb_4 c57 (.A(net938),
    .B(net29),
    .C_N(net30),
    .D_N(net17),
    .X(net32));
 sky130_fd_sc_hd__and3b_4 c570 (.A_N(net536),
    .B(net804),
    .C(net859),
    .X(net545));
 sky130_fd_sc_hd__or3_2 c571 (.A(net112),
    .B(net545),
    .C(net859),
    .X(net546));
 sky130_fd_sc_hd__or3b_1 c572 (.A(clknet_1_0__leaf_net426),
    .B(net986),
    .C_N(net249),
    .X(net547));
 sky130_fd_sc_hd__nor3_1 c573 (.A(net518),
    .B(net400),
    .C(net999),
    .Y(net548));
 sky130_fd_sc_hd__and3b_4 c574 (.A_N(net543),
    .B(clknet_1_0__leaf_net547),
    .C(net788),
    .X(net549));
 sky130_fd_sc_hd__and3b_4 c575 (.A_N(net545),
    .B(clknet_1_1__leaf_net426),
    .C(clknet_1_0__leaf_net431),
    .X(net550));
 sky130_fd_sc_hd__buf_2 c576 (.A(net896),
    .X(net551));
 sky130_fd_sc_hd__or4bb_2 c577 (.A(clknet_1_1__leaf_net435),
    .B(net413),
    .C_N(net538),
    .D_N(clknet_1_0__leaf_net547),
    .X(net552));
 sky130_fd_sc_hd__nor3_4 c578 (.A(clknet_1_1__leaf_net531),
    .B(net551),
    .C(net420),
    .Y(net553));
 sky130_fd_sc_hd__or3_1 c579 (.A(net543),
    .B(net125),
    .C(net986),
    .X(net554));
 sky130_fd_sc_hd__or4bb_2 c58 (.A(net26),
    .B(net27),
    .C_N(net23),
    .D_N(net25),
    .X(net33));
 sky130_fd_sc_hd__mux4_4 c580 (.A0(net298),
    .A1(clknet_1_1__leaf_net431),
    .A2(net420),
    .A3(net551),
    .S0(clknet_1_0__leaf_net547),
    .S1(net543),
    .X(net555));
 sky130_fd_sc_hd__nand3b_1 c581 (.A_N(net986),
    .B(net133),
    .C(net999),
    .Y(net556));
 sky130_fd_sc_hd__or4bb_2 c582 (.A(net1000),
    .B(net551),
    .C_N(clknet_1_0__leaf_net435),
    .D_N(net803),
    .X(net557));
 sky130_fd_sc_hd__nor3_2 c583 (.A(net420),
    .B(clknet_1_1__leaf_net557),
    .C(clknet_1_1__leaf_net426),
    .Y(net558));
 sky130_fd_sc_hd__sdfbbn_2 c584 (.CLK_N(clknet_4_6_0_clk),
    .D(net551),
    .RESET_B(net948),
    .SCD(clknet_1_0__leaf_net558),
    .SCE(clknet_1_0__leaf_net547),
    .SET_B(net796),
    .Q(net560),
    .Q_N(net559));
 sky130_fd_sc_hd__mux4_2 c585 (.A0(clknet_1_1__leaf_net435),
    .A1(net545),
    .A2(clknet_1_1__leaf_net557),
    .A3(net551),
    .S0(net559),
    .S1(net858),
    .X(net561));
 sky130_fd_sc_hd__or3_1 c586 (.A(net26),
    .B(net554),
    .C(clknet_1_1__leaf_net513),
    .X(net562));
 sky130_fd_sc_hd__or4bb_4 c587 (.A(clknet_1_0__leaf_net562),
    .B(net552),
    .C_N(clknet_1_1__leaf_net557),
    .D_N(clknet_1_0__leaf_net547),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_1 c588 (.A(net896),
    .X(net564));
 sky130_fd_sc_hd__or3b_2 c589 (.A(clknet_1_0__leaf_net557),
    .B(net134),
    .C_N(clknet_1_1__leaf_net513),
    .X(net565));
 sky130_fd_sc_hd__a2111o_1 c59 (.A1(net28),
    .A2(net23),
    .B1(net11),
    .C1(net24),
    .D1(net27),
    .X(net34));
 sky130_fd_sc_hd__sdfstp_2 c590 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net562),
    .SCD(clknet_1_1__leaf_net557),
    .SCE(net26),
    .SET_B(net1015),
    .Q(net566));
 sky130_fd_sc_hd__mux4_2 c591 (.A0(net256),
    .A1(net564),
    .A2(net298),
    .A3(clknet_1_0__leaf_net549),
    .S0(clknet_1_0__leaf_net557),
    .S1(net831),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 c592 (.A(net903),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net523),
    .A1(net568),
    .A2(net401),
    .A3(net566),
    .S0(net420),
    .S1(clknet_1_1__leaf_net860),
    .X(net569));
 sky130_fd_sc_hd__sdfstp_4 c594 (.CLK(clknet_4_6_0_clk),
    .D(net556),
    .SCD(net560),
    .SCE(clknet_1_0__leaf_net565),
    .SET_B(net1014),
    .Q(net570));
 sky130_fd_sc_hd__and3_1 c595 (.A(net174),
    .B(net452),
    .C(net413),
    .X(net571));
 sky130_fd_sc_hd__or3_1 c596 (.A(net532),
    .B(net979),
    .C(net566),
    .X(net957));
 sky130_fd_sc_hd__sdfbbn_1 c597 (.CLK_N(clknet_4_6_0_clk),
    .D(net556),
    .RESET_B(clknet_1_1__leaf_net529),
    .SCD(net452),
    .SCE(net545),
    .SET_B(net412),
    .Q(net573),
    .Q_N(net572));
 sky130_fd_sc_hd__or4bb_1 c598 (.A(net135),
    .B(net386),
    .C_N(net413),
    .D_N(net786),
    .X(net574));
 sky130_fd_sc_hd__or4bb_4 c599 (.A(net530),
    .B(net412),
    .C_N(net176),
    .D_N(net125),
    .X(net575));
 sky130_fd_sc_hd__or4bb_4 c60 (.A(net23),
    .B(net29),
    .C_N(net34),
    .D_N(net5),
    .X(net35));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(clknet_1_1__leaf_net171),
    .A1(net570),
    .A2(net1029),
    .A3(net575),
    .S0(net997),
    .S1(net999),
    .X(net576));
 sky130_fd_sc_hd__or4bb_4 c601 (.A(net176),
    .B(net444),
    .C_N(clknet_1_1__leaf_net171),
    .D_N(net451),
    .X(net577));
 sky130_fd_sc_hd__or4bb_2 c602 (.A(net412),
    .B(net13),
    .C_N(clknet_1_0__leaf_net576),
    .D_N(net193),
    .X(net578));
 sky130_fd_sc_hd__sedfxbp_2 c603 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_0__leaf_net576),
    .DE(net175),
    .SCD(net997),
    .SCE(net1028),
    .Q(net580),
    .Q_N(net579));
 sky130_fd_sc_hd__sedfxbp_1 c604 (.CLK(clknet_4_6_0_clk),
    .D(net401),
    .DE(net979),
    .SCD(clknet_1_0__leaf_net565),
    .SCE(net786),
    .Q(net582),
    .Q_N(net581));
 sky130_fd_sc_hd__or4bb_1 c605 (.A(net574),
    .B(net579),
    .C_N(net801),
    .D_N(net835),
    .X(net583));
 sky130_fd_sc_hd__or4bb_1 c606 (.A(net193),
    .B(net13),
    .C_N(net579),
    .D_N(net840),
    .X(net584));
 sky130_fd_sc_hd__o2111ai_1 c607 (.A1(net254),
    .A2(net573),
    .B1(clknet_1_1__leaf_net171),
    .C1(clknet_1_1__leaf_net576),
    .D1(clknet_1_1__leaf_net842),
    .Y(net585));
 sky130_fd_sc_hd__mux4_4 c608 (.A0(net583),
    .A1(net580),
    .A2(net984),
    .A3(net575),
    .S0(net572),
    .S1(clknet_1_0__leaf_net842),
    .X(net586));
 sky130_fd_sc_hd__a2111o_2 c609 (.A1(net577),
    .A2(net115),
    .B1(net574),
    .C1(clknet_1_0__leaf_net586),
    .D1(net979),
    .X(net587));
 sky130_fd_sc_hd__or4bb_1 c61 (.A(net35),
    .B(net34),
    .C_N(net26),
    .D_N(net25),
    .X(net36));
 sky130_fd_sc_hd__sedfxtp_1 c610 (.CLK(clknet_4_6_0_clk),
    .D(net413),
    .DE(clknet_1_0__leaf_net587),
    .SCD(clknet_1_1__leaf_net576),
    .SCE(net999),
    .Q(net588));
 sky130_fd_sc_hd__a2111o_2 c611 (.A1(net573),
    .A2(net1021),
    .B1(net538),
    .C1(clknet_1_1__leaf_net576),
    .D1(clknet_1_0__leaf_net586),
    .X(net589));
 sky130_fd_sc_hd__sdfbbp_1 c612 (.CLK(clknet_4_6_0_clk),
    .D(net1020),
    .RESET_B(clknet_1_1__leaf_net589),
    .SCD(net580),
    .SCE(clknet_1_1__leaf_net586),
    .SET_B(clknet_1_0__leaf_net585),
    .Q(net590));
 sky130_fd_sc_hd__sdfbbn_1 c613 (.CLK_N(clknet_4_6_0_clk),
    .D(net588),
    .RESET_B(clknet_1_0__leaf_net587),
    .SCD(net581),
    .SCE(clknet_1_0__leaf_net589),
    .SET_B(net254),
    .Q(net591));
 sky130_fd_sc_hd__sedfxtp_1 c614 (.CLK(clknet_4_6_0_clk),
    .D(net511),
    .DE(net591),
    .SCD(clknet_1_1__leaf_net587),
    .SCE(clknet_1_0__leaf_net586),
    .Q(net592));
 sky130_fd_sc_hd__or4bb_4 c615 (.A(net14),
    .B(net590),
    .C_N(net560),
    .D_N(clknet_1_0__leaf_net446),
    .X(net593));
 sky130_fd_sc_hd__a2111oi_2 c616 (.A1(net461),
    .A2(net204),
    .B1(clknet_1_0__leaf_net593),
    .C1(net473),
    .D1(clknet_1_0__leaf_net958),
    .Y(net594));
 sky130_fd_sc_hd__a2111o_4 c617 (.A1(net571),
    .A2(clknet_1_1__leaf_net594),
    .B1(net948),
    .C1(net559),
    .D1(net831),
    .X(net595));
 sky130_fd_sc_hd__or4bb_4 c618 (.A(clknet_1_0__leaf_net463),
    .B(clknet_1_0__leaf_net593),
    .C_N(net834),
    .D_N(clknet_1_1__leaf_net844),
    .X(net596));
 sky130_fd_sc_hd__a2111oi_2 c619 (.A1(net282),
    .A2(net79),
    .B1(clknet_1_1__leaf_net596),
    .C1(net461),
    .D1(net831),
    .Y(net597));
 sky130_fd_sc_hd__a2111o_1 c62 (.A1(net34),
    .A2(net31),
    .B1(net36),
    .C1(net27),
    .D1(net21),
    .X(net37));
 sky130_fd_sc_hd__sedfxtp_1 c620 (.CLK(clknet_4_6_0_clk),
    .D(net175),
    .DE(clknet_1_0__leaf_net594),
    .SCD(clknet_1_0__leaf_net595),
    .SCE(net249),
    .Q(net598));
 sky130_fd_sc_hd__sdfrbp_1 c621 (.CLK(clknet_4_13_0_clk),
    .D(clknet_1_0__leaf_net558),
    .RESET_B(net282),
    .SCD(clknet_1_1__leaf_net553),
    .SCE(net204),
    .Q(net600),
    .Q_N(net599));
 sky130_fd_sc_hd__mux4_4 c622 (.A0(net597),
    .A1(clknet_1_0__leaf_net561),
    .A2(clknet_1_0__leaf_net553),
    .A3(clknet_1_1__leaf_net529),
    .S0(net282),
    .S1(clknet_1_1__leaf_net844),
    .X(net601));
 sky130_fd_sc_hd__o2111ai_2 c623 (.A1(net249),
    .A2(clknet_1_0__leaf_net553),
    .B1(net570),
    .C1(net598),
    .D1(net801),
    .Y(net951));
 sky130_fd_sc_hd__o2111ai_4 c624 (.A1(net560),
    .A2(clknet_1_0__leaf_net596),
    .B1(clknet_1_0__leaf_net951),
    .C1(net449),
    .D1(net570),
    .Y(net602));
 sky130_fd_sc_hd__a2111o_1 c625 (.A1(clknet_1_1__leaf_net553),
    .A2(net592),
    .B1(clknet_1_0__leaf_net463),
    .C1(net599),
    .D1(clknet_1_0__leaf_net951),
    .X(net603));
 sky130_fd_sc_hd__a2111oi_0 c626 (.A1(net249),
    .A2(clknet_1_0__leaf_net951),
    .B1(clknet_1_1__leaf_net558),
    .C1(net948),
    .D1(net826),
    .Y(net604));
 sky130_fd_sc_hd__sdfbbn_1 c627 (.CLK_N(clknet_4_15_0_clk),
    .D(net54),
    .RESET_B(net175),
    .SCD(clknet_1_1__leaf_net593),
    .SCE(clknet_1_1__leaf_net844),
    .SET_B(net849),
    .Q(net969));
 sky130_fd_sc_hd__o2111a_4 c628 (.A1(net461),
    .A2(clknet_1_0__leaf_net951),
    .B1(clknet_1_0__leaf_net958),
    .C1(clknet_1_1__leaf_net844),
    .D1(net850),
    .X(net605));
 sky130_fd_sc_hd__sdfbbp_1 c629 (.CLK(clknet_4_13_0_clk),
    .D(clknet_1_1__leaf_net561),
    .RESET_B(net922),
    .SCD(clknet_1_0__leaf_net603),
    .SCE(net79),
    .SET_B(net1016),
    .Q(net607),
    .Q_N(net606));
 sky130_fd_sc_hd__a2111oi_1 c63 (.A1(net17),
    .A2(net33),
    .B1(net35),
    .C1(net22),
    .D1(net798),
    .Y(net38));
 sky130_fd_sc_hd__mux4_2 c630 (.A0(clknet_1_1__leaf_net602),
    .A1(clknet_1_0__leaf_net951),
    .A2(net559),
    .A3(net606),
    .S0(net789),
    .S1(net831),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net204),
    .A1(net339),
    .A2(net474),
    .A3(net321),
    .S0(net606),
    .S1(clknet_1_1__leaf_net951),
    .X(net947));
 sky130_fd_sc_hd__a2111oi_4 c632 (.A1(net79),
    .A2(clknet_1_0__leaf_net605),
    .B1(net204),
    .C1(net606),
    .D1(net790),
    .Y(net609));
 sky130_fd_sc_hd__mux4_4 c633 (.A0(net600),
    .A1(clknet_1_1__leaf_net595),
    .A2(net339),
    .A3(clknet_1_1__leaf_net609),
    .S0(clknet_1_0__leaf_net608),
    .S1(clknet_1_1__leaf_net605),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(clknet_1_0__leaf_net608),
    .A1(clknet_1_0__leaf_net609),
    .A2(net606),
    .A3(net204),
    .S0(clknet_1_0__leaf_net958),
    .S1(net831),
    .X(net954));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net598),
    .A1(clknet_1_0__leaf_net602),
    .A2(clknet_1_0__leaf_net463),
    .A3(clknet_1_0__leaf_net951),
    .S0(clknet_1_0__leaf_net609),
    .S1(clknet_1_0__leaf_net605),
    .X(net611));
 sky130_fd_sc_hd__o2111ai_4 c636 (.A1(clknet_1_1__leaf_net609),
    .A2(net610),
    .B1(clknet_1_1__leaf_net608),
    .C1(clknet_1_1__leaf_net951),
    .D1(clknet_1_1__leaf_net605),
    .Y(net612));
 sky130_fd_sc_hd__a2111oi_1 c637 (.A1(clknet_1_1__leaf_net603),
    .A2(clknet_1_1__leaf_net605),
    .B1(clknet_1_0__leaf_net947),
    .C1(clknet_1_0__leaf_net612),
    .D1(clknet_1_1__leaf_net609),
    .Y(net613));
 sky130_fd_sc_hd__mux4_1 c64 (.A0(net972),
    .A1(net34),
    .A2(net24),
    .A3(net12),
    .S0(net35),
    .X(net39));
 sky130_fd_sc_hd__or2b_4 c65 (.A(net943),
    .B_N(net17),
    .X(net40));
 sky130_fd_sc_hd__or2_2 c66 (.A(net25),
    .B(net988),
    .X(net41));
 sky130_fd_sc_hd__nand2_2 c660 (.A(net382),
    .B(clknet_1_0__leaf_net513),
    .Y(net614));
 sky130_fd_sc_hd__nand2_1 c661 (.A(net118),
    .B(net857),
    .Y(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 c662 (.A(net805),
    .X(net616));
 sky130_fd_sc_hd__and3_1 c663 (.A(net512),
    .B(net616),
    .C(net253),
    .X(net617));
 sky130_fd_sc_hd__nand2_1 c664 (.A(net253),
    .B(net984),
    .Y(net618));
 sky130_fd_sc_hd__buf_16 c665 (.A(net805),
    .X(net619));
 sky130_fd_sc_hd__or2b_1 c666 (.A(net944),
    .B_N(net512),
    .X(net620));
 sky130_fd_sc_hd__and3_1 c667 (.A(net114),
    .B(net619),
    .C(clknet_1_0__leaf_net513),
    .X(net621));
 sky130_fd_sc_hd__buf_8 c668 (.A(clknet_1_0__leaf_net756),
    .X(net622));
 sky130_fd_sc_hd__or2_2 c669 (.A(net253),
    .B(net382),
    .X(net623));
 sky130_fd_sc_hd__and2b_1 c67 (.A_N(net50),
    .B(net937),
    .X(net42));
 sky130_fd_sc_hd__or2_2 c670 (.A(net507),
    .B(net617),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__nand3b_1 c672 (.A_N(clknet_1_0__leaf_net622),
    .B(net125),
    .C(net624),
    .Y(net626));
 sky130_fd_sc_hd__or2b_1 c673 (.A(net1013),
    .B_N(net512),
    .X(net627));
 sky130_fd_sc_hd__or2b_1 c674 (.A(net616),
    .B_N(net624),
    .X(net628));
 sky130_fd_sc_hd__nand3_2 c675 (.A(net617),
    .B(net616),
    .C(net857),
    .Y(net629));
 sky130_fd_sc_hd__or3_2 c676 (.A(net627),
    .B(net386),
    .C(net616),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd1_1 c677 (.A(clknet_1_0__leaf_net919),
    .X(net631));
 sky130_fd_sc_hd__buf_6 c678 (.A(net813),
    .X(net632));
 sky130_fd_sc_hd__mux4_2 c679 (.A0(net522),
    .A1(clknet_1_1__leaf_net622),
    .A2(clknet_1_0__leaf_net631),
    .A3(clknet_1_1__leaf_net519),
    .S0(net624),
    .S1(net379),
    .X(net633));
 sky130_fd_sc_hd__or2_1 c68 (.A(net58),
    .B(net11),
    .X(net43));
 sky130_fd_sc_hd__or3b_1 c680 (.A(clknet_1_0__leaf_net630),
    .B(net617),
    .C_N(net805),
    .X(net634));
 sky130_fd_sc_hd__inv_12 c671_13 (.A(clknet_1_1__leaf_net756),
    .Y(net1013));
 sky130_fd_sc_hd__buf_1 c682 (.A(net743),
    .X(net636));
 sky130_fd_sc_hd__nand3b_2 c683 (.A_N(net654),
    .B(net632),
    .C(clknet_1_1__leaf_net862),
    .Y(net637));
 sky130_fd_sc_hd__a2111oi_1 c684 (.A1(net624),
    .A2(net546),
    .B1(net993),
    .C1(net858),
    .D1(clknet_1_0__leaf_net862),
    .Y(net638));
 sky130_fd_sc_hd__clkbuf_1 c685 (.A(net916),
    .X(net639));
 sky130_fd_sc_hd__nor3b_4 c686 (.A(net656),
    .B(clknet_1_0__leaf_net634),
    .C_N(net857),
    .Y(net640));
 sky130_fd_sc_hd__sdfrbp_1 c687 (.CLK(clknet_4_5_0_clk),
    .D(net639),
    .RESET_B(net618),
    .SCD(clknet_1_0__leaf_net640),
    .SCE(net993),
    .Q(net642),
    .Q_N(net641));
 sky130_fd_sc_hd__buf_4 c688 (.A(net813),
    .X(net643));
 sky130_fd_sc_hd__or4bb_4 c689 (.A(clknet_1_1__leaf_net640),
    .B(net654),
    .C_N(net656),
    .D_N(net993),
    .X(net644));
 sky130_fd_sc_hd__nand2_1 c69 (.A(net59),
    .B(net61),
    .Y(net44));
 sky130_fd_sc_hd__or4bb_4 c690 (.A(net619),
    .B(clknet_1_1__leaf_net655),
    .C_N(net654),
    .D_N(net534),
    .X(net645));
 sky130_fd_sc_hd__inv_6 c691 (.A(net916),
    .Y(net646));
 sky130_fd_sc_hd__clkbuf_1 c692 (.A(net913),
    .X(net647));
 sky130_fd_sc_hd__inv_2 c693 (.A(net906),
    .Y(net648));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(clknet_1_0__leaf_net655),
    .A1(net646),
    .A2(net642),
    .A3(clknet_1_1__leaf_net638),
    .S0(clknet_1_0__leaf_net544),
    .S1(net993),
    .X(net649));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net647),
    .A1(net147),
    .A2(net646),
    .A3(net619),
    .S0(net993),
    .S1(net813),
    .X(net650));
 sky130_fd_sc_hd__buf_2 c696 (.A(net744),
    .X(net651));
 sky130_fd_sc_hd__or3b_1 c697 (.A(net936),
    .B(net537),
    .C_N(net619),
    .X(net652));
 sky130_fd_sc_hd__or3b_4 c698 (.A(net624),
    .B(net993),
    .C_N(net833),
    .X(net653));
 sky130_fd_sc_hd__nor3b_2 c699 (.A(net534),
    .B(net14),
    .C_N(net993),
    .Y(net654));
 sky130_fd_sc_hd__inv_4 c70 (.A(net794),
    .Y(net45));
 sky130_fd_sc_hd__or4bb_2 c700 (.A(net521),
    .B(net1012),
    .C_N(net632),
    .D_N(clknet_1_0__leaf_net513),
    .X(net655));
 sky130_fd_sc_hd__inv_4 c701 (.A(net914),
    .Y(net656));
 sky130_fd_sc_hd__buf_6 c702 (.A(net909),
    .X(net657));
 sky130_fd_sc_hd__mux4_4 c703 (.A0(net618),
    .A1(net654),
    .A2(net125),
    .A3(clknet_1_0__leaf_net529),
    .S0(net993),
    .S1(net858),
    .X(net658));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net537),
    .A1(clknet_1_0__leaf_net550),
    .A2(net392),
    .A3(net657),
    .S0(clknet_1_0__leaf_net547),
    .S1(net636),
    .X(net659));
 sky130_fd_sc_hd__a2111o_4 c705 (.A1(net636),
    .A2(clknet_1_1__leaf_net547),
    .B1(clknet_1_1__leaf_net634),
    .C1(net981),
    .D1(net857),
    .X(net660));
 sky130_fd_sc_hd__a2111oi_1 c706 (.A1(net292),
    .A2(net551),
    .B1(net648),
    .C1(net994),
    .D1(net629),
    .Y(net661));
 sky130_fd_sc_hd__sdfbbn_1 c707 (.CLK_N(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net621),
    .RESET_B(clknet_1_0__leaf_net544),
    .SCD(net392),
    .SCE(net857),
    .SET_B(clknet_1_0__leaf_net861),
    .Q(net663),
    .Q_N(net662));
 sky130_fd_sc_hd__a2111o_1 c708 (.A1(clknet_1_1__leaf_net513),
    .A2(net643),
    .B1(net651),
    .C1(net994),
    .D1(net857),
    .X(net664));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net392),
    .A1(net651),
    .A2(net1011),
    .A3(net40),
    .S0(net995),
    .S1(clknet_1_0__leaf_net547),
    .X(net665));
 sky130_fd_sc_hd__and2_1 c71 (.A(net42),
    .B(net798),
    .X(net46));
 sky130_fd_sc_hd__sdfbbn_1 c710 (.CLK_N(clknet_4_5_0_clk),
    .D(net296),
    .RESET_B(clknet_1_1__leaf_net634),
    .SCD(clknet_1_1__leaf_net664),
    .SCE(net386),
    .SET_B(net994),
    .Q(net667),
    .Q_N(net666));
 sky130_fd_sc_hd__sdfbbp_1 c711 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net664),
    .RESET_B(net661),
    .SCD(net386),
    .SCE(net651),
    .SET_B(net786),
    .Q(net669),
    .Q_N(net668));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net40),
    .A1(net657),
    .A2(net537),
    .A3(net668),
    .S0(net653),
    .S1(net566),
    .X(net670));
 sky130_fd_sc_hd__sdfbbn_1 c713 (.CLK_N(clknet_4_5_0_clk),
    .D(net665),
    .RESET_B(net147),
    .SCD(net1023),
    .SCE(net999),
    .SET_B(net857),
    .Q(net672),
    .Q_N(net671));
 sky130_fd_sc_hd__o2111ai_4 c714 (.A1(net1010),
    .A2(net569),
    .B1(net667),
    .C1(net296),
    .D1(net648),
    .Y(net673));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net629),
    .A1(net981),
    .A2(net672),
    .A3(net643),
    .S0(clknet_1_0__leaf_net664),
    .S1(clknet_1_0__leaf_net673),
    .X(net674));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net629),
    .A1(net546),
    .A2(net40),
    .A3(clknet_1_1__leaf_net637),
    .S0(clknet_1_0__leaf_net673),
    .S1(net778),
    .X(net675));
 sky130_fd_sc_hd__mux4_4 c717 (.A0(net672),
    .A1(clknet_1_1__leaf_net673),
    .A2(clknet_1_0__leaf_net529),
    .A3(clknet_1_1__leaf_net634),
    .S0(net994),
    .S1(net857),
    .X(net676));
 sky130_fd_sc_hd__a2111oi_2 c718 (.A1(net546),
    .A2(clknet_1_0__leaf_net673),
    .B1(net551),
    .C1(net643),
    .D1(net657),
    .Y(net677));
 sky130_fd_sc_hd__mux4_2 c719 (.A0(net653),
    .A1(net632),
    .A2(clknet_1_0__leaf_net673),
    .A3(net993),
    .S0(net785),
    .S1(net864),
    .X(net678));
 sky130_fd_sc_hd__and2b_1 c72 (.A_N(net11),
    .B(net45),
    .X(net47));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net669),
    .A1(clknet_1_1__leaf_net565),
    .A2(net994),
    .A3(clknet_1_1__leaf_net673),
    .S0(clknet_1_0__leaf_net677),
    .S1(net866),
    .X(net679));
 sky130_fd_sc_hd__mux4_4 c721 (.A0(net978),
    .A1(clknet_1_0__leaf_net673),
    .A2(clknet_1_0__leaf_net547),
    .A3(net671),
    .S0(net648),
    .S1(net785),
    .X(net680));
 sky130_fd_sc_hd__mux4_2 c722 (.A0(net653),
    .A1(clknet_1_1__leaf_net565),
    .A2(clknet_1_0__leaf_net673),
    .A3(net566),
    .S0(net777),
    .S1(net857),
    .X(net681));
 sky130_fd_sc_hd__mux4_4 c723 (.A0(net680),
    .A1(clknet_1_1__leaf_net550),
    .A2(clknet_1_0__leaf_net634),
    .A3(net657),
    .S0(clknet_1_0__leaf_net673),
    .S1(net863),
    .X(net682));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net632),
    .A1(clknet_1_1__leaf_net673),
    .A2(net666),
    .A3(clknet_1_0__leaf_net547),
    .S0(net867),
    .S1(net869),
    .X(net683));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net683),
    .A1(clknet_1_1__leaf_net673),
    .A2(net971),
    .A3(net865),
    .S0(net868),
    .S1(net869),
    .X(net684));
 sky130_fd_sc_hd__a2111oi_2 c726 (.A1(net452),
    .A2(clknet_1_0__leaf_net565),
    .B1(net449),
    .C1(net971),
    .D1(net545),
    .Y(net685));
 sky130_fd_sc_hd__mux4_2 c727 (.A0(net386),
    .A1(net984),
    .A2(clknet_1_0__leaf_net659),
    .A3(net942),
    .S0(net997),
    .S1(net575),
    .X(net686));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(clknet_1_1__leaf_net677),
    .A1(net971),
    .A2(net575),
    .A3(clknet_1_1__leaf_net446),
    .S0(net785),
    .S1(net870),
    .X(net687));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(clknet_1_0__leaf_net659),
    .A1(net580),
    .A2(clknet_1_0__leaf_net565),
    .A3(net575),
    .S0(clknet_1_1__leaf_net547),
    .S1(net994),
    .X(net688));
 sky130_fd_sc_hd__or2_1 c73 (.A(net47),
    .B(net46),
    .X(net48));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_1__leaf_net637),
    .A1(net16),
    .A2(clknet_1_1__leaf_net446),
    .A3(net984),
    .S0(net451),
    .S1(net870),
    .X(net689));
 sky130_fd_sc_hd__o2111a_1 c731 (.A1(net643),
    .A2(net997),
    .B1(net545),
    .C1(net994),
    .D1(net871),
    .X(net690));
 sky130_fd_sc_hd__sdfbbn_1 c732 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net586),
    .RESET_B(net545),
    .SCD(net984),
    .SCE(net570),
    .SET_B(net971),
    .Q(net692),
    .Q_N(net691));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net575),
    .A1(net663),
    .A2(net971),
    .A3(net994),
    .S0(net984),
    .S1(clknet_1_1__leaf_net544),
    .X(net693));
 sky130_fd_sc_hd__a2111oi_2 c734 (.A1(net566),
    .A2(clknet_1_0__leaf_net446),
    .B1(net579),
    .C1(net871),
    .D1(net875),
    .Y(net694));
 sky130_fd_sc_hd__mux4_4 c735 (.A0(net9),
    .A1(net971),
    .A2(clknet_1_0__leaf_net694),
    .A3(net566),
    .S0(net994),
    .S1(net871),
    .X(net695));
 sky130_fd_sc_hd__mux4_2 c736 (.A0(clknet_1_1__leaf_net585),
    .A1(net971),
    .A2(net691),
    .A3(net514),
    .S0(net871),
    .S1(net876),
    .X(net696));
 sky130_fd_sc_hd__mux4_2 c737 (.A0(net995),
    .A1(net575),
    .A2(clknet_1_1__leaf_net659),
    .A3(clknet_1_1__leaf_net586),
    .S0(net877),
    .S1(net878),
    .X(net697));
 sky130_fd_sc_hd__sdfbbp_1 c738 (.CLK(clknet_4_7_0_clk),
    .D(net514),
    .RESET_B(net9),
    .SCD(clknet_1_0__leaf_net694),
    .SCE(net971),
    .SET_B(net1017),
    .Q(net699),
    .Q_N(net698));
 sky130_fd_sc_hd__mux4_2 c739 (.A0(net667),
    .A1(net514),
    .A2(net623),
    .A3(clknet_1_0__leaf_net808),
    .S0(net874),
    .S1(net878),
    .X(net700));
 sky130_fd_sc_hd__inv_1 c74 (.A(net793),
    .Y(net49));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net699),
    .A1(net579),
    .A2(net995),
    .A3(net870),
    .S0(net871),
    .S1(net878),
    .X(net701));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net648),
    .A1(clknet_1_1__leaf_net547),
    .A2(net698),
    .A3(net871),
    .S0(net878),
    .S1(net879),
    .X(net702));
 sky130_fd_sc_hd__sdfbbn_1 c742 (.CLK_N(clknet_4_7_0_clk),
    .D(net660),
    .RESET_B(net699),
    .SCD(clknet_1_0__leaf_net702),
    .SCE(clknet_1_1__leaf_net808),
    .SET_B(net878),
    .Q(net703));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net580),
    .A1(net663),
    .A2(net994),
    .A3(clknet_1_0__leaf_net702),
    .S0(net878),
    .S1(net880),
    .X(net704));
 sky130_fd_sc_hd__mux4_4 c744 (.A0(net703),
    .A1(clknet_1_1__leaf_net702),
    .A2(net451),
    .A3(net691),
    .S0(net666),
    .S1(net876),
    .X(net705));
 sky130_fd_sc_hd__mux4_4 c745 (.A0(net690),
    .A1(clknet_1_1__leaf_net544),
    .A2(clknet_1_0__leaf_net702),
    .A3(net623),
    .S0(net871),
    .S1(net883),
    .X(net706));
 sky130_fd_sc_hd__mux4_2 c746 (.A0(net701),
    .A1(clknet_1_1__leaf_net446),
    .A2(clknet_1_1__leaf_net702),
    .A3(net878),
    .S0(net883),
    .S1(net884),
    .X(net707));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_1__leaf_net446),
    .A1(net662),
    .A2(clknet_1_1__leaf_net702),
    .A3(net881),
    .S0(net882),
    .S1(net885),
    .X(net708));
 sky130_fd_sc_hd__mux4_2 c748 (.A0(net692),
    .A1(clknet_1_0__leaf_net612),
    .A2(net16),
    .A3(clknet_1_1__leaf_net198),
    .S0(net473),
    .S1(net872),
    .X(net709));
 sky130_fd_sc_hd__mux4_2 c749 (.A0(net339),
    .A1(net458),
    .A2(net613),
    .A3(clknet_1_1__leaf_net198),
    .S0(net570),
    .S1(net941),
    .X(net710));
 sky130_fd_sc_hd__or2_4 c75 (.A(net45),
    .B(net55),
    .X(net946));
 sky130_fd_sc_hd__mux4_2 c750 (.A0(net607),
    .A1(clknet_1_1__leaf_net612),
    .A2(net570),
    .A3(net834),
    .S0(net873),
    .S1(net886),
    .X(net711));
 sky130_fd_sc_hd__mux4_4 c751 (.A0(net709),
    .A1(clknet_1_1__leaf_net694),
    .A2(clknet_1_1__leaf_net198),
    .A3(net105),
    .S0(net809),
    .S1(clknet_1_1__leaf_net861),
    .X(net712));
 sky130_fd_sc_hd__mux4_2 c752 (.A0(net474),
    .A1(net651),
    .A2(net942),
    .A3(net997),
    .S0(clknet_1_0__leaf_net861),
    .S1(net887),
    .X(net713));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net611),
    .A1(net474),
    .A2(net785),
    .A3(clknet_1_1__leaf_net861),
    .S0(net869),
    .S1(net887),
    .X(net714));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net713),
    .A1(net474),
    .A2(net607),
    .A3(net786),
    .S0(net873),
    .S1(net887),
    .X(net715));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net922),
    .A1(clknet_1_1__leaf_net547),
    .A2(clknet_1_1__leaf_net529),
    .A3(net826),
    .S0(net871),
    .S1(net887),
    .X(net716));
 sky130_fd_sc_hd__mux4_4 c756 (.A0(net711),
    .A1(net570),
    .A2(net997),
    .A3(clknet_1_1__leaf_net529),
    .S0(clknet_1_1__leaf_net547),
    .S1(net888),
    .X(net717));
 sky130_fd_sc_hd__mux4_4 c757 (.A0(net570),
    .A1(net115),
    .A2(net715),
    .A3(clknet_1_1__leaf_net694),
    .S0(net886),
    .S1(net887),
    .X(net718));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net607),
    .A1(clknet_1_1__leaf_net718),
    .A2(clknet_1_1__leaf_net547),
    .A3(net570),
    .S0(net887),
    .S1(net889),
    .X(net719));
 sky130_fd_sc_hd__mux4_4 c759 (.A0(clknet_1_1__leaf_net529),
    .A1(net449),
    .A2(clknet_1_0__leaf_net718),
    .A3(net570),
    .S0(net887),
    .S1(net889),
    .X(net720));
 sky130_fd_sc_hd__or2_2 c76 (.A(net930),
    .B(net22),
    .X(net50));
 sky130_fd_sc_hd__mux4_4 c760 (.A0(net321),
    .A1(net714),
    .A2(net692),
    .A3(clknet_1_0__leaf_net718),
    .S0(net889),
    .S1(net890),
    .X(net721));
 sky130_fd_sc_hd__mux4_4 c761 (.A0(net657),
    .A1(clknet_1_1__leaf_net547),
    .A2(net719),
    .A3(net607),
    .S0(clknet_1_1__leaf_net718),
    .S1(net889),
    .X(net722));
 sky130_fd_sc_hd__mux4_2 c762 (.A0(net721),
    .A1(clknet_1_1__leaf_net198),
    .A2(clknet_1_1__leaf_net529),
    .A3(net939),
    .S0(net889),
    .S1(net891),
    .X(net723));
 sky130_fd_sc_hd__nand2b_1 c77 (.A_N(net14),
    .B(net41),
    .Y(net51));
 sky130_fd_sc_hd__clkbuf_1 c78 (.A(net794),
    .X(net52));
 sky130_fd_sc_hd__and2b_1 c79 (.A_N(net41),
    .B(net19),
    .X(net53));
 sky130_fd_sc_hd__nor2_2 c80 (.A(net932),
    .B(net928),
    .Y(net54));
 sky130_fd_sc_hd__nor2_1 c81 (.A(net942),
    .B(net22),
    .Y(net55));
 sky130_fd_sc_hd__nor3_1 c82 (.A(net53),
    .B(net51),
    .C(net937),
    .Y(net56));
 sky130_fd_sc_hd__and2b_1 c83 (.A_N(net53),
    .B(net932),
    .X(net57));
 sky130_fd_sc_hd__and2_1 c84 (.A(net57),
    .B(net798),
    .X(net58));
 sky130_fd_sc_hd__and2b_1 c85 (.A_N(net51),
    .B(net57),
    .X(net59));
 sky130_fd_sc_hd__and2b_1 c86 (.A_N(net55),
    .B(net59),
    .X(net60));
 sky130_fd_sc_hd__inv_1 c87 (.A(net751),
    .Y(net61));
 sky130_fd_sc_hd__or2b_1 c88 (.A(net46),
    .B_N(net798),
    .X(net62));
 sky130_fd_sc_hd__inv_4 c89 (.A(net814),
    .Y(net63));
 sky130_fd_sc_hd__or2_2 c90 (.A(net926),
    .B(net46),
    .X(net64));
 sky130_fd_sc_hd__nor2_1 c91 (.A(net62),
    .B(net64),
    .Y(net65));
 sky130_fd_sc_hd__and2_1 c92 (.A(net65),
    .B(net63),
    .X(net66));
 sky130_fd_sc_hd__nor2b_1 c93 (.A(net33),
    .B_N(net934),
    .Y(net67));
 sky130_fd_sc_hd__nand2b_2 c94 (.A_N(net63),
    .B(net926),
    .Y(net68));
 sky130_fd_sc_hd__nor2_1 c95 (.A(net17),
    .B(net68),
    .Y(net69));
 sky130_fd_sc_hd__or2_1 c96 (.A(net64),
    .B(net62),
    .X(net70));
 sky130_fd_sc_hd__nand2_1 c97 (.A(net922),
    .B(net798),
    .Y(net71));
 sky130_fd_sc_hd__and2b_1 c98 (.A_N(net65),
    .B(net68),
    .X(net72));
 sky130_fd_sc_hd__and2b_1 c99 (.A_N(net64),
    .B(net68),
    .X(net73));
 sky130_fd_sc_hd__mux4_4 merge763 (.A0(net30),
    .A1(net220),
    .A2(clknet_1_0__leaf_net233),
    .A3(clknet_1_0__leaf_net358),
    .S0(net308),
    .S1(net821),
    .X(net724));
 sky130_fd_sc_hd__mux4_4 merge764 (.A0(net1003),
    .A1(net101),
    .A2(net220),
    .A3(net191),
    .S0(net237),
    .S1(net226),
    .X(net725));
 sky130_fd_sc_hd__sdfrtn_1 merge765 (.CLK_N(clknet_4_8_0_clk),
    .D(net177),
    .RESET_B(net43),
    .SCD(net151),
    .SCE(clknet_1_0__leaf_net213),
    .Q(net726));
 sky130_fd_sc_hd__sdfbbn_1 merge766 (.CLK_N(clknet_4_9_0_clk),
    .D(net217),
    .RESET_B(net332),
    .SCD(net83),
    .SCE(net333),
    .SET_B(net1025),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__or4bb_2 merge767 (.A(net311),
    .B(net147),
    .C_N(net315),
    .D_N(clknet_1_1__leaf_net168),
    .X(net729));
 sky130_fd_sc_hd__mux4_2 merge768 (.A0(net328),
    .A1(net179),
    .A2(net979),
    .A3(clknet_1_1__leaf_net167),
    .S0(net118),
    .S1(net183),
    .X(net730));
 sky130_fd_sc_hd__sdfrtp_1 merge769 (.CLK(clknet_4_2_0_clk),
    .D(net152),
    .RESET_B(clknet_1_0__leaf_net167),
    .SCD(net143),
    .SCE(net179),
    .Q(net731));
 sky130_fd_sc_hd__sdfrtp_1 merge770 (.CLK(clknet_4_8_0_clk),
    .D(net77),
    .RESET_B(net69),
    .SCD(net90),
    .SCE(net89),
    .Q(net732));
 sky130_fd_sc_hd__or4bb_2 merge771 (.A(net379),
    .B(net518),
    .C_N(net387),
    .D_N(clknet_1_0__leaf_net529),
    .X(net733));
 sky130_fd_sc_hd__or3b_1 merge772 (.A(clknet_1_0__leaf_net519),
    .B(net114),
    .C_N(net615),
    .X(net734));
 sky130_fd_sc_hd__or4bb_1 merge773 (.A(net303),
    .B(net308),
    .C_N(net289),
    .D_N(clknet_1_0__leaf_net295),
    .X(net735));
 sky130_fd_sc_hd__mux4_2 merge774 (.A0(clknet_1_0__leaf_net431),
    .A1(net298),
    .A2(net518),
    .A3(clknet_1_1__leaf_net549),
    .S0(clknet_1_0__leaf_net557),
    .S1(net795),
    .X(net736));
 sky130_fd_sc_hd__or4bb_1 merge775 (.A(net43),
    .B(net35),
    .C_N(net11),
    .D_N(net1031),
    .X(net737));
 sky130_fd_sc_hd__mux4_2 merge776 (.A0(net393),
    .A1(net148),
    .A2(net135),
    .A3(net397),
    .S0(clknet_1_0__leaf_net395),
    .S1(net378),
    .X(net738));
 sky130_fd_sc_hd__mux4_1 merge777 (.A0(net934),
    .A1(net379),
    .A2(net1000),
    .A3(net516),
    .S0(net383),
    .S1(net807),
    .X(net739));
 sky130_fd_sc_hd__mux4_4 merge778 (.A0(net152),
    .A1(net7),
    .A2(net155),
    .A3(net150),
    .S0(net14),
    .S1(net147),
    .X(net740));
 sky130_fd_sc_hd__or4bb_1 merge779 (.A(net381),
    .B(net118),
    .C_N(net377),
    .D_N(net383),
    .X(net741));
 sky130_fd_sc_hd__mux4_1 merge780 (.A0(net271),
    .A1(net146),
    .A2(net991),
    .A3(net283),
    .S0(net123),
    .S1(net112),
    .X(net742));
 sky130_fd_sc_hd__sdfbbp_1 merge781 (.CLK(clknet_4_4_0_clk),
    .D(net971),
    .RESET_B(clknet_1_0__leaf_net621),
    .SCD(net4),
    .SCE(net545),
    .SET_B(net653),
    .Q(net744),
    .Q_N(net743));
 sky130_fd_sc_hd__or4bb_4 merge782 (.A(net166),
    .B(net256),
    .C_N(clknet_1_1__leaf_net389),
    .D_N(clknet_1_1__leaf_net390),
    .X(net745));
 sky130_fd_sc_hd__sdfrtp_4 merge783 (.CLK(clknet_4_2_0_clk),
    .D(net291),
    .RESET_B(net290),
    .SCD(net275),
    .SCE(net146),
    .Q(net746));
 sky130_fd_sc_hd__sdfsbp_1 merge784 (.CLK(clknet_4_2_0_clk),
    .D(net27),
    .SCD(clknet_1_0__leaf_net168),
    .SCE(net419),
    .SET_B(net287),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__sdfsbp_1 merge785 (.CLK(clknet_4_1_0_clk),
    .D(net528),
    .SCD(net959),
    .SCE(net935),
    .SET_B(net535),
    .Q(net750),
    .Q_N(net749));
 sky130_fd_sc_hd__sdfstp_1 merge786 (.CLK(clknet_4_8_0_clk),
    .D(net89),
    .SCD(net64),
    .SCE(net60),
    .SET_B(net926),
    .Q(net751));
 sky130_fd_sc_hd__mux4_4 merge787 (.A0(net127),
    .A1(clknet_1_0__leaf_net529),
    .A2(net383),
    .A3(net262),
    .S0(net379),
    .S1(net833),
    .X(net752));
 sky130_fd_sc_hd__mux4_1 merge788 (.A0(net51),
    .A1(clknet_1_0__leaf_net430),
    .A2(net989),
    .A3(net195),
    .S0(net249),
    .S1(clknet_1_1__leaf_net390),
    .X(net753));
 sky130_fd_sc_hd__or4bb_1 merge789 (.A(net974),
    .B(net936),
    .C_N(net91),
    .D_N(net93),
    .X(net754));
 sky130_fd_sc_hd__or4bb_1 merge790 (.A(net56),
    .B(net44),
    .C_N(net48),
    .D_N(net328),
    .X(net755));
 sky130_fd_sc_hd__dlymetal6s2s_1 merge791 (.A(clknet_1_0__leaf_net920),
    .X(net756));
 sky130_fd_sc_hd__mux4_2 merge792 (.A0(net566),
    .A1(clknet_1_0__leaf_net565),
    .A2(net304),
    .A3(net280),
    .S0(net254),
    .S1(clknet_1_0__leaf_net860),
    .X(net757));
 sky130_fd_sc_hd__mux4_2 merge793 (.A0(net286),
    .A1(net394),
    .A2(clknet_1_1__leaf_net395),
    .A3(net290),
    .S0(net19),
    .S1(net306),
    .X(net758));
 sky130_fd_sc_hd__mux4_1 merge794 (.A0(net533),
    .A1(net528),
    .A2(net949),
    .A3(net646),
    .S0(clknet_1_0__leaf_net637),
    .S1(net782),
    .X(net759));
 sky130_fd_sc_hd__mux4_4 merge795 (.A0(net319),
    .A1(clknet_1_0__leaf_net295),
    .A2(net183),
    .A3(net247),
    .S0(net996),
    .S1(net535),
    .X(net760));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(net318),
    .A1(net998),
    .A2(net309),
    .A3(net336),
    .S0(clknet_1_0__leaf_net341),
    .S1(net340),
    .X(net761));
 sky130_fd_sc_hd__mux4_2 merge797 (.A0(net535),
    .A1(net534),
    .A2(net533),
    .A3(net147),
    .S0(net386),
    .S1(clknet_1_1__leaf_net513),
    .X(net762));
 sky130_fd_sc_hd__mux4_2 merge798 (.A0(net210),
    .A1(clknet_1_0__leaf_net208),
    .A2(net214),
    .A3(net200),
    .S0(net30),
    .S1(net137),
    .X(net763));
 sky130_fd_sc_hd__mux4_4 merge799 (.A0(net63),
    .A1(net926),
    .A2(net32),
    .A3(net98),
    .S0(net94),
    .S1(net162),
    .X(net764));
 sky130_fd_sc_hd__mux4_1 merge800 (.A0(net628),
    .A1(net993),
    .A2(clknet_1_1__leaf_net640),
    .A3(net643),
    .S0(net782),
    .S1(net833),
    .X(net765));
 sky130_fd_sc_hd__sdfbbn_1 merge801 (.CLK_N(clknet_4_12_0_clk),
    .D(net447),
    .RESET_B(net946),
    .SCD(net1029),
    .SCE(net974),
    .SET_B(net193),
    .Q(net767),
    .Q_N(net766));
 sky130_fd_sc_hd__mux4_4 merge802 (.A0(clknet_1_1__leaf_net168),
    .A1(net41),
    .A2(clknet_1_0__leaf_net295),
    .A3(net164),
    .S0(net183),
    .S1(net173),
    .X(net768));
 sky130_fd_sc_hd__mux4_4 merge803 (.A0(net654),
    .A1(net656),
    .A2(net653),
    .A3(net641),
    .S0(net651),
    .S1(clknet_1_0__leaf_net637),
    .X(net769));
 sky130_fd_sc_hd__mux4_2 merge804 (.A0(net526),
    .A1(net535),
    .A2(net316),
    .A3(net987),
    .S0(clknet_1_0__leaf_net295),
    .S1(net779),
    .X(net770));
 sky130_fd_sc_hd__mux4_2 merge805 (.A0(net314),
    .A1(net316),
    .A2(net998),
    .A3(net96),
    .S0(net955),
    .S1(net100),
    .X(net771));
 sky130_fd_sc_hd__mux4_4 merge806 (.A0(net614),
    .A1(clknet_1_1__leaf_net631),
    .A2(clknet_1_1__leaf_net630),
    .A3(clknet_1_0__leaf_net638),
    .S0(net545),
    .S1(clknet_1_0__leaf_net640),
    .X(net772));
 sky130_fd_sc_hd__mux4_4 merge807 (.A0(net259),
    .A1(net971),
    .A2(clknet_1_0__leaf_net621),
    .A3(net975),
    .S0(net532),
    .S1(net535),
    .X(net773));
 sky130_fd_sc_hd__mux4_1 merge808 (.A0(net626),
    .A1(net624),
    .A2(clknet_1_0__leaf_net634),
    .A3(net379),
    .S0(net521),
    .S1(net620),
    .X(net774));
 sky130_fd_sc_hd__dfrbp_1 merge809 (.CLK(clknet_4_2_0_clk),
    .D(net169),
    .Q(net172),
    .Q_N(net775));
 sky130_fd_sc_hd__dfrbp_1 merge810 (.CLK(clknet_4_5_0_clk),
    .D(net670),
    .RESET_B(net674),
    .Q(net778),
    .Q_N(net777));
 sky130_fd_sc_hd__dfrtn_1 merge811 (.CLK_N(clknet_4_1_0_clk),
    .D(net540),
    .RESET_B(net733),
    .Q(net779));
 sky130_fd_sc_hd__dfrtp_1 merge812 (.CLK(clknet_4_14_0_clk),
    .D(net467),
    .RESET_B(net477),
    .Q(net780));
 sky130_fd_sc_hd__dfrtp_1 merge813 (.CLK(clknet_4_2_0_clk),
    .D(net437),
    .Q(net443));
 sky130_fd_sc_hd__dfrtp_1 merge814 (.CLK(clknet_4_5_0_clk),
    .D(net644),
    .RESET_B(net645),
    .Q(net782));
 sky130_fd_sc_hd__dfsbp_1 merge815 (.CLK(clknet_4_2_0_clk),
    .D(net735),
    .SET_B(net745),
    .Q(net784),
    .Q_N(net783));
 sky130_fd_sc_hd__dfsbp_2 merge816 (.CLK(clknet_4_3_0_clk),
    .D(net424),
    .SET_B(net436),
    .Q(net786),
    .Q_N(net785));
 sky130_fd_sc_hd__dfstp_1 merge817 (.CLK(clknet_4_11_0_clk),
    .D(net503),
    .SET_B(net488),
    .Q(net968));
 sky130_fd_sc_hd__dfstp_1 merge818 (.CLK(clknet_4_10_0_clk),
    .D(net97),
    .SET_B(net104),
    .Q(net787));
 sky130_fd_sc_hd__dfstp_1 merge819 (.CLK(clknet_4_1_0_clk),
    .D(net525),
    .SET_B(net739),
    .Q(net788));
 sky130_fd_sc_hd__dlrbn_1 merge820 (.D(net601),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net604),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__dlrbn_1 merge821 (.D(net194),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net189),
    .Q(net792),
    .Q_N(net791));
 sky130_fd_sc_hd__dlrbp_2 merge822 (.D(net737),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net755),
    .Q(net794),
    .Q_N(net793));
 sky130_fd_sc_hd__dlrbp_1 merge823 (.D(net555),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net563),
    .Q(net796),
    .Q_N(net795));
 sky130_fd_sc_hd__dlrtn_1 merge824 (.D(net322),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net729),
    .Q(net797));
 sky130_fd_sc_hd__dlrtn_1 merge825 (.D(net37),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net39));
 sky130_fd_sc_hd__dlrtn_1 merge826 (.D(net343),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net346),
    .Q(net799));
 sky130_fd_sc_hd__dlrtp_1 merge827 (.D(net209),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net212),
    .Q(net800));
 sky130_fd_sc_hd__dlrtp_1 merge828 (.D(net578),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net584),
    .Q(net801));
 sky130_fd_sc_hd__dlrtp_1 merge829 (.D(net228),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net234),
    .Q(net802));
 sky130_fd_sc_hd__edfxbp_1 merge830 (.CLK(clknet_4_1_0_clk),
    .D(net406),
    .DE(net407),
    .Q(net804),
    .Q_N(net803));
 sky130_fd_sc_hd__edfxtp_1 merge831 (.CLK(clknet_4_4_0_clk),
    .D(net633),
    .DE(net734),
    .Q(net805));
 sky130_fd_sc_hd__sdlclkp_1 merge832 (.CLK(clknet_4_11_0_clk),
    .GATE(net363),
    .SCE(net364),
    .GCLK(net806));
 sky130_fd_sc_hd__sdlclkp_2 merge833 (.CLK(clknet_4_1_0_clk),
    .GATE(net385),
    .GCLK(net391));
 sky130_fd_sc_hd__sdlclkp_4 merge834 (.CLK(clknet_4_6_0_clk),
    .GATE(net685),
    .SCE(net688),
    .GCLK(net808));
 sky130_fd_sc_hd__dfrbp_1 merge835 (.CLK(clknet_4_15_0_clk),
    .D(net723),
    .RESET_B(net710),
    .Q(net809));
 sky130_fd_sc_hd__dfrbp_2 merge836 (.CLK(clknet_4_0_0_clk),
    .D(net741),
    .RESET_B(net742),
    .Q(net811),
    .Q_N(net810));
 sky130_fd_sc_hd__dfrtn_1 merge837 (.CLK_N(clknet_4_11_0_clk),
    .D(net454),
    .RESET_B(net497),
    .Q(net812));
 sky130_fd_sc_hd__dfrtp_1 merge838 (.CLK(clknet_4_5_0_clk),
    .D(net649),
    .RESET_B(net772),
    .Q(net813));
 sky130_fd_sc_hd__dfrtp_4 merge839 (.CLK(clknet_4_8_0_clk),
    .D(net218),
    .RESET_B(net754),
    .Q(net814));
 sky130_fd_sc_hd__dfrtp_1 merge840 (.CLK(clknet_4_0_0_clk),
    .D(net411),
    .Q(net414));
 sky130_fd_sc_hd__dfxbp_1 s841 (.CLK(clknet_4_10_0_clk),
    .D(net102),
    .Q(net817),
    .Q_N(net816));
 sky130_fd_sc_hd__dfxbp_1 s842 (.CLK(clknet_4_10_0_clk),
    .D(net103),
    .Q(net819),
    .Q_N(net818));
 sky130_fd_sc_hd__dfxtp_1 s843 (.CLK(clknet_4_2_0_clk),
    .D(net188),
    .Q(net820));
 sky130_fd_sc_hd__dfxtp_2 s844 (.CLK(clknet_4_11_0_clk),
    .D(net330),
    .Q(net821));
 sky130_fd_sc_hd__dfxtp_1 s845 (.CLK(clknet_4_9_0_clk),
    .D(net348),
    .Q(net822));
 sky130_fd_sc_hd__dlclkp_1 s846 (.CLK(clknet_4_9_0_clk),
    .GATE(net349),
    .GCLK(net823));
 sky130_fd_sc_hd__dlclkp_2 s847 (.CLK(clknet_4_11_0_clk),
    .GATE(net350),
    .GCLK(net958));
 sky130_fd_sc_hd__dlclkp_4 s848 (.CLK(clknet_4_11_0_clk),
    .GATE(net351),
    .GCLK(net824));
 sky130_fd_sc_hd__dlxbn_1 s849 (.D(net352),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net826),
    .Q_N(net825));
 sky130_fd_sc_hd__dlxbn_1 s850 (.D(net365),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net828),
    .Q_N(net827));
 sky130_fd_sc_hd__dlxbp_1 s851 (.D(net368),
    .GATE(clknet_4_11_0_clk),
    .Q(net829));
 sky130_fd_sc_hd__dlxtn_1 s852 (.D(net370),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net830));
 sky130_fd_sc_hd__dlxtn_4 s853 (.D(net408),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net831));
 sky130_fd_sc_hd__dlxtn_1 s854 (.D(net409),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net832));
 sky130_fd_sc_hd__dlxtp_1 s855 (.D(net410),
    .GATE(clknet_4_1_0_clk),
    .Q(net833));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s856 (.D(net434),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net834));
 sky130_fd_sc_hd__dfxbp_1 s857 (.CLK(clknet_4_3_0_clk),
    .D(net441),
    .Q(net836),
    .Q_N(net835));
 sky130_fd_sc_hd__dfxbp_1 s858 (.CLK(clknet_4_3_0_clk),
    .D(net453),
    .Q(net838),
    .Q_N(net837));
 sky130_fd_sc_hd__dfxtp_1 s859 (.CLK(clknet_4_3_0_clk),
    .D(net455),
    .Q(net839));
 sky130_fd_sc_hd__dfxtp_1 s860 (.CLK(clknet_4_12_0_clk),
    .D(net456),
    .Q(net840));
 sky130_fd_sc_hd__dfxtp_1 s861 (.CLK(clknet_4_12_0_clk),
    .D(net457),
    .Q(net841));
 sky130_fd_sc_hd__dlclkp_1 s862 (.CLK(clknet_4_3_0_clk),
    .GATE(net459),
    .GCLK(net842));
 sky130_fd_sc_hd__dlclkp_2 s863 (.CLK(clknet_4_14_0_clk),
    .GATE(net464),
    .GCLK(net843));
 sky130_fd_sc_hd__dlclkp_4 s864 (.CLK(clknet_4_14_0_clk),
    .GATE(net471),
    .GCLK(net844));
 sky130_fd_sc_hd__dlxbn_1 s865 (.D(net483),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net846),
    .Q_N(net845));
 sky130_fd_sc_hd__dlxbn_1 s866 (.D(net485),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net848),
    .Q_N(net847));
 sky130_fd_sc_hd__dlxbp_1 s867 (.D(net487),
    .GATE(clknet_4_15_0_clk),
    .Q(net850),
    .Q_N(net849));
 sky130_fd_sc_hd__dlxtn_1 s868 (.D(net490),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net851));
 sky130_fd_sc_hd__dlxtn_1 s869 (.D(net491),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net852));
 sky130_fd_sc_hd__dlxtn_1 s870 (.D(net492),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net853));
 sky130_fd_sc_hd__dlxtp_1 s871 (.D(net495),
    .GATE(clknet_4_11_0_clk),
    .Q(net960));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s872 (.D(net496),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net854));
 sky130_fd_sc_hd__dfxbp_1 s873 (.CLK(clknet_4_11_0_clk),
    .D(net501),
    .Q(net964),
    .Q_N(net855));
 sky130_fd_sc_hd__dfxbp_1 s874 (.CLK(clknet_4_11_0_clk),
    .D(net502),
    .Q(net952),
    .Q_N(net856));
 sky130_fd_sc_hd__dfxtp_4 s875 (.CLK(clknet_4_4_0_clk),
    .D(net524),
    .Q(net857));
 sky130_fd_sc_hd__dfxtp_1 s876 (.CLK(clknet_4_4_0_clk),
    .D(net541),
    .Q(net858));
 sky130_fd_sc_hd__dfxtp_1 s877 (.CLK(clknet_4_1_0_clk),
    .D(net542),
    .Q(net859));
 sky130_fd_sc_hd__dlclkp_1 s878 (.CLK(clknet_4_3_0_clk),
    .GATE(net567),
    .GCLK(net860));
 sky130_fd_sc_hd__dlclkp_2 s879 (.CLK(clknet_4_5_0_clk),
    .GATE(net650),
    .GCLK(net861));
 sky130_fd_sc_hd__dlclkp_4 s880 (.CLK(clknet_4_4_0_clk),
    .GATE(net658),
    .GCLK(net862));
 sky130_fd_sc_hd__dlxbn_1 s881 (.D(net675),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net864),
    .Q_N(net863));
 sky130_fd_sc_hd__dlxbn_1 s882 (.D(net676),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net865));
 sky130_fd_sc_hd__dlxbp_1 s883 (.D(net678),
    .GATE(clknet_4_5_0_clk),
    .Q(net866));
 sky130_fd_sc_hd__dlxtn_1 s884 (.D(net679),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net867));
 sky130_fd_sc_hd__dlxtn_1 s885 (.D(net681),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net868));
 sky130_fd_sc_hd__dlxtn_1 s886 (.D(net682),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net869));
 sky130_fd_sc_hd__dlxtp_1 s887 (.D(net684),
    .GATE(clknet_4_7_0_clk),
    .Q(net870));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s888 (.D(net686),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net871));
 sky130_fd_sc_hd__dfxbp_1 s889 (.CLK(clknet_4_13_0_clk),
    .D(net687),
    .Q(net873),
    .Q_N(net872));
 sky130_fd_sc_hd__dfxbp_1 s890 (.CLK(clknet_4_7_0_clk),
    .D(net689),
    .Q(net875),
    .Q_N(net874));
 sky130_fd_sc_hd__dfxtp_1 s891 (.CLK(clknet_4_7_0_clk),
    .D(net693),
    .Q(net876));
 sky130_fd_sc_hd__dfxtp_1 s892 (.CLK(clknet_4_7_0_clk),
    .D(net695),
    .Q(net877));
 sky130_fd_sc_hd__dfxtp_2 s893 (.CLK(clknet_4_7_0_clk),
    .D(net696),
    .Q(net878));
 sky130_fd_sc_hd__dlclkp_1 s894 (.CLK(clknet_4_7_0_clk),
    .GATE(net697),
    .GCLK(net879));
 sky130_fd_sc_hd__dlclkp_2 s895 (.CLK(clknet_4_7_0_clk),
    .GATE(net700),
    .GCLK(net880));
 sky130_fd_sc_hd__dlclkp_4 s896 (.CLK(clknet_4_13_0_clk),
    .GATE(net704),
    .GCLK(net881));
 sky130_fd_sc_hd__dlxbn_1 s897 (.D(net705),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net883),
    .Q_N(net882));
 sky130_fd_sc_hd__dlxbn_1 s898 (.D(net706),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net884));
 sky130_fd_sc_hd__dlxbp_1 s899 (.D(net707),
    .GATE(clknet_4_7_0_clk),
    .Q(net885));
 sky130_fd_sc_hd__dlxtn_1 s900 (.D(net708),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net886));
 sky130_fd_sc_hd__dlxtn_2 s901 (.D(net712),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net887));
 sky130_fd_sc_hd__dlxtn_1 s902 (.D(net716),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net888));
 sky130_fd_sc_hd__dlxtp_1 s903 (.D(net717),
    .GATE(clknet_4_15_0_clk),
    .Q(net889));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s904 (.D(net720),
    .SLEEP_B(clknet_4_15_0_clk),
    .Q(net890));
 sky130_fd_sc_hd__dfxbp_1 s905 (.CLK(clknet_4_15_0_clk),
    .D(net722),
    .Q(net891));
 sky130_fd_sc_hd__dfxbp_1 s906 (.CLK(clknet_4_10_0_clk),
    .D(net724),
    .Q(net893),
    .Q_N(net892));
 sky130_fd_sc_hd__dfxtp_1 s907 (.CLK(clknet_4_10_0_clk),
    .D(net725),
    .Q(net894));
 sky130_fd_sc_hd__dfxtp_2 s908 (.CLK(clknet_4_12_0_clk),
    .D(net730),
    .Q(net895));
 sky130_fd_sc_hd__dfxtp_1 s909 (.CLK(clknet_4_4_0_clk),
    .D(net736),
    .Q(net896));
 sky130_fd_sc_hd__dlclkp_1 s910 (.CLK(clknet_4_0_0_clk),
    .GATE(net738),
    .GCLK(net897));
 sky130_fd_sc_hd__dlclkp_2 s911 (.CLK(clknet_4_2_0_clk),
    .GATE(net740),
    .GCLK(net898));
 sky130_fd_sc_hd__dlclkp_4 s912 (.CLK(clknet_4_1_0_clk),
    .GATE(net752),
    .GCLK(net899));
 sky130_fd_sc_hd__dlxbn_1 s913 (.D(net753),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net901),
    .Q_N(net900));
 sky130_fd_sc_hd__dlxbn_1 s914 (.D(net757),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net903),
    .Q_N(net902));
 sky130_fd_sc_hd__dlxbp_1 s915 (.D(net758),
    .GATE(clknet_4_0_0_clk),
    .Q(net905),
    .Q_N(net904));
 sky130_fd_sc_hd__dlxtn_1 s916 (.D(net759),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net906));
 sky130_fd_sc_hd__dlxtn_1 s917 (.D(net760),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net907));
 sky130_fd_sc_hd__dlxtn_1 s918 (.D(net761),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net908));
 sky130_fd_sc_hd__dlxtp_1 s919 (.D(net762),
    .GATE(clknet_4_4_0_clk),
    .Q(net909));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s920 (.D(net763),
    .SLEEP_B(clknet_4_8_0_clk),
    .Q(net910));
 sky130_fd_sc_hd__dfxbp_1 s921 (.CLK(clknet_4_10_0_clk),
    .D(net764),
    .Q(net912),
    .Q_N(net911));
 sky130_fd_sc_hd__dfxbp_1 s922 (.CLK(clknet_4_5_0_clk),
    .D(net765),
    .Q(net914),
    .Q_N(net913));
 sky130_fd_sc_hd__dfxtp_1 s923 (.CLK(clknet_4_9_0_clk),
    .D(net768),
    .Q(net915));
 sky130_fd_sc_hd__dfxtp_1 s924 (.CLK(clknet_4_5_0_clk),
    .D(net769),
    .Q(net916));
 sky130_fd_sc_hd__dfxtp_2 s925 (.CLK(clknet_4_0_0_clk),
    .D(net770),
    .Q(net917));
 sky130_fd_sc_hd__dlclkp_1 s926 (.CLK(clknet_4_8_0_clk),
    .GATE(net771),
    .GCLK(net918));
 sky130_fd_sc_hd__dlclkp_2 s927 (.CLK(clknet_4_4_0_clk),
    .GATE(net773),
    .GCLK(net919));
 sky130_fd_sc_hd__dlclkp_4 s928 (.CLK(clknet_4_4_0_clk),
    .GATE(net774),
    .GCLK(net920));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(in0),
    .X(net921));
 sky130_fd_sc_hd__buf_4 input2 (.A(in1),
    .X(net922));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net923));
 sky130_fd_sc_hd__buf_1 input4 (.A(in11),
    .X(net924));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net925));
 sky130_fd_sc_hd__buf_2 input6 (.A(in13),
    .X(net926));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(in14),
    .X(net927));
 sky130_fd_sc_hd__buf_4 input8 (.A(in15),
    .X(net928));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(in16),
    .X(net929));
 sky130_fd_sc_hd__buf_2 input10 (.A(in17),
    .X(net930));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net931));
 sky130_fd_sc_hd__buf_4 input12 (.A(in19),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(in2),
    .X(net933));
 sky130_fd_sc_hd__buf_2 input14 (.A(in20),
    .X(net934));
 sky130_fd_sc_hd__buf_2 input15 (.A(in21),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_8 input16 (.A(in22),
    .X(net936));
 sky130_fd_sc_hd__buf_2 input17 (.A(in23),
    .X(net937));
 sky130_fd_sc_hd__buf_1 input18 (.A(in24),
    .X(net938));
 sky130_fd_sc_hd__buf_4 input19 (.A(in3),
    .X(net939));
 sky130_fd_sc_hd__buf_1 input20 (.A(in4),
    .X(net940));
 sky130_fd_sc_hd__buf_4 input21 (.A(in5),
    .X(net941));
 sky130_fd_sc_hd__buf_4 input22 (.A(in6),
    .X(net942));
 sky130_fd_sc_hd__buf_4 input23 (.A(in7),
    .X(net943));
 sky130_fd_sc_hd__buf_2 input24 (.A(in8),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in9),
    .X(net945));
 sky130_fd_sc_hd__buf_2 output26 (.A(net946),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(clknet_1_1__leaf_net947),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output28 (.A(net990),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output29 (.A(net949),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(clknet_1_1__leaf_net950),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(clknet_1_1__leaf_net951),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output32 (.A(net952),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output33 (.A(net953),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net954),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output35 (.A(net955),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(clknet_1_1__leaf_net956),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output37 (.A(net957),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(clknet_1_1__leaf_net958),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output39 (.A(net959),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output40 (.A(net960),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output41 (.A(net961),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output42 (.A(net962),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net963),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output44 (.A(net964),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output45 (.A(net965),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(clknet_1_1__leaf_net966),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net967),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output48 (.A(net968),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output49 (.A(net969),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(clknet_1_1__leaf_net970),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net623),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_1 wire52 (.A(net973),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_1 max_cap53 (.A(net38),
    .X(net973));
 sky130_fd_sc_hd__buf_4 fanout54 (.A(net32),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_1 max_cap55 (.A(net1032),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_2 max_cap56 (.A(net450),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_2 max_cap57 (.A(net146),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_1 max_cap58 (.A(net1033),
    .X(net978));
 sky130_fd_sc_hd__buf_4 fanout59 (.A(net282),
    .X(net979));
 sky130_fd_sc_hd__buf_1 wire60 (.A(net281),
    .X(net980));
 sky130_fd_sc_hd__buf_1 wire61 (.A(net548),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_2 max_cap62 (.A(net279),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net371),
    .X(net983));
 sky130_fd_sc_hd__buf_4 fanout64 (.A(net514),
    .X(net984));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(net203),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_2 max_cap66 (.A(net265),
    .X(net986));
 sky130_fd_sc_hd__buf_2 fanout67 (.A(net153),
    .X(net987));
 sky130_fd_sc_hd__buf_4 fanout68 (.A(net16),
    .X(net988));
 sky130_fd_sc_hd__buf_4 fanout69 (.A(net248),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(net948),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(net270),
    .X(net991));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(net131),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_4 fanout73 (.A(net995),
    .X(net993));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(net995),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(net652),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_2 max_cap76 (.A(net413),
    .X(net996));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(net321),
    .X(net997));
 sky130_fd_sc_hd__buf_2 fanout78 (.A(net320),
    .X(net998));
 sky130_fd_sc_hd__buf_4 fanout79 (.A(net834),
    .X(net999));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(net105),
    .X(net1000));
 sky130_fd_sc_hd__clkinv_8 c180_1 (.A(clknet_1_0__leaf_net898),
    .Y(net1001));
 sky130_fd_sc_hd__clkinv_8 net999_2 (.A(clknet_1_0__leaf_net898),
    .Y(net1002));
 sky130_fd_sc_hd__clkinv_16 c187_4 (.A(clknet_1_1__leaf_net898),
    .Y(net1004));
 sky130_fd_sc_hd__clkinv_16 c187_5 (.A(clknet_1_0__leaf_net898),
    .Y(net1005));
 sky130_fd_sc_hd__clkinv_16 c187_6 (.A(clknet_1_0__leaf_net898),
    .Y(net1006));
 sky130_fd_sc_hd__clkinv_16 c187_7 (.A(clknet_1_0__leaf_net898),
    .Y(net1007));
 sky130_fd_sc_hd__inv_1 c344_9 (.A(net918),
    .Y(net1009));
 sky130_fd_sc_hd__clkinv_1 c681_11 (.A(clknet_1_1__leaf_net920),
    .Y(net1011));
 sky130_fd_sc_hd__clkinv_1 c681_12 (.A(clknet_1_0__leaf_net920),
    .Y(net1012));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net920 (.A(net920),
    .X(clknet_0_net920));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net920 (.A(clknet_0_net920),
    .X(clknet_1_0__leaf_net920));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net920 (.A(clknet_0_net920),
    .X(clknet_1_1__leaf_net920));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net655 (.A(net655),
    .X(clknet_0_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net673 (.A(net673),
    .X(clknet_0_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_0__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net673 (.A(clknet_0_net673),
    .X(clknet_1_1__leaf_net673));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net677 (.A(net677),
    .X(clknet_0_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_0__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_1__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net756 (.A(net756),
    .X(clknet_0_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net756 (.A(clknet_0_net756),
    .X(clknet_1_0__leaf_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net756 (.A(clknet_0_net756),
    .X(clknet_1_1__leaf_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net630 (.A(net630),
    .X(clknet_0_net630));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net630 (.A(clknet_0_net630),
    .X(clknet_1_0__leaf_net630));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net630 (.A(clknet_0_net630),
    .X(clknet_1_1__leaf_net630));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net634 (.A(net634),
    .X(clknet_0_net634));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net634 (.A(clknet_0_net634),
    .X(clknet_1_0__leaf_net634));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net634 (.A(clknet_0_net634),
    .X(clknet_1_1__leaf_net634));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net640 (.A(net640),
    .X(clknet_0_net640));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net640 (.A(clknet_0_net640),
    .X(clknet_1_0__leaf_net640));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net640 (.A(clknet_0_net640),
    .X(clknet_1_1__leaf_net640));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net622 (.A(net622),
    .X(clknet_0_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_0__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_1__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net919 (.A(net919),
    .X(clknet_0_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net919 (.A(clknet_0_net919),
    .X(clknet_1_0__leaf_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net919 (.A(clknet_0_net919),
    .X(clknet_1_1__leaf_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net631 (.A(net631),
    .X(clknet_0_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net631 (.A(clknet_0_net631),
    .X(clknet_1_0__leaf_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net631 (.A(clknet_0_net631),
    .X(clknet_1_1__leaf_net631));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net544 (.A(net544),
    .X(clknet_0_net544));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net544 (.A(clknet_0_net544),
    .X(clknet_1_0__leaf_net544));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net544 (.A(clknet_0_net544),
    .X(clknet_1_1__leaf_net544));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net324 (.A(net324),
    .X(clknet_0_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net324 (.A(clknet_0_net324),
    .X(clknet_1_0__leaf_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net324 (.A(clknet_0_net324),
    .X(clknet_1_1__leaf_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net475 (.A(net475),
    .X(clknet_0_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net475 (.A(clknet_0_net475),
    .X(clknet_1_0__leaf_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net475 (.A(clknet_0_net475),
    .X(clknet_1_1__leaf_net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net843 (.A(net843),
    .X(clknet_0_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net843 (.A(clknet_0_net843),
    .X(clknet_1_0__leaf_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net843 (.A(clknet_0_net843),
    .X(clknet_1_1__leaf_net843));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net472 (.A(net472),
    .X(clknet_0_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_0__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_1__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net956 (.A(net956),
    .X(clknet_0_net956));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net956 (.A(clknet_0_net956),
    .X(clknet_1_0__leaf_net956));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net956 (.A(clknet_0_net956),
    .X(clknet_1_1__leaf_net956));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net478 (.A(net478),
    .X(clknet_0_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_0__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_1__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net476 (.A(net476),
    .X(clknet_0_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net476 (.A(clknet_0_net476),
    .X(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net476 (.A(clknet_0_net476),
    .X(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net327 (.A(net327),
    .X(clknet_0_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net531 (.A(net531),
    .X(clknet_0_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net531 (.A(clknet_0_net531),
    .X(clknet_1_0__leaf_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net531 (.A(clknet_0_net531),
    .X(clknet_1_1__leaf_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net553 (.A(net553),
    .X(clknet_0_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_0__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_1__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net603 (.A(net603),
    .X(clknet_0_net603));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net603 (.A(clknet_0_net603),
    .X(clknet_1_0__leaf_net603));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net603 (.A(clknet_0_net603),
    .X(clknet_1_1__leaf_net603));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net951 (.A(net951),
    .X(clknet_0_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net951 (.A(clknet_0_net951),
    .X(clknet_1_0__leaf_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net951 (.A(clknet_0_net951),
    .X(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net612 (.A(net612),
    .X(clknet_0_net612));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net612 (.A(clknet_0_net612),
    .X(clknet_1_0__leaf_net612));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net612 (.A(clknet_0_net612),
    .X(clknet_1_1__leaf_net612));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net947 (.A(net947),
    .X(clknet_0_net947));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net947 (.A(clknet_0_net947),
    .X(clknet_1_0__leaf_net947));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net947 (.A(clknet_0_net947),
    .X(clknet_1_1__leaf_net947));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net608 (.A(net608),
    .X(clknet_0_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net608 (.A(clknet_0_net608),
    .X(clknet_1_0__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net608 (.A(net625),
    .X(clknet_1_1__leaf_net608));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net605 (.A(net605),
    .X(clknet_0_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_0__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_1__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net609 (.A(net609),
    .X(clknet_0_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_0__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_1__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net602 (.A(net602),
    .X(clknet_0_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net602 (.A(net323),
    .X(clknet_1_0__leaf_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net602 (.A(clknet_0_net602),
    .X(clknet_1_1__leaf_net602));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net388 (.A(net388),
    .X(clknet_0_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net388 (.A(clknet_0_net388),
    .X(clknet_1_0__leaf_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net388 (.A(clknet_0_net388),
    .X(clknet_1_1__leaf_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net508 (.A(net508),
    .X(clknet_0_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_0__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_1__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net519 (.A(net519),
    .X(clknet_0_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_1__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net513 (.A(net513),
    .X(clknet_0_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_0__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_1__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net664 (.A(net664),
    .X(clknet_0_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_0__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_1__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net621 (.A(net621),
    .X(clknet_0_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net621 (.A(clknet_0_net621),
    .X(clknet_1_0__leaf_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net621 (.A(clknet_0_net621),
    .X(clknet_1_1__leaf_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net565 (.A(net565),
    .X(clknet_0_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net565 (.A(clknet_0_net565),
    .X(clknet_1_0__leaf_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net565 (.A(clknet_0_net565),
    .X(clknet_1_1__leaf_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net808 (.A(net808),
    .X(clknet_0_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net808 (.A(clknet_0_net808),
    .X(clknet_1_0__leaf_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net808 (.A(clknet_0_net808),
    .X(clknet_1_1__leaf_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net529 (.A(net529),
    .X(clknet_0_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net529 (.A(clknet_0_net529),
    .X(clknet_1_0__leaf_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net529 (.A(clknet_0_net529),
    .X(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net862 (.A(net862),
    .X(clknet_0_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net862 (.A(clknet_0_net862),
    .X(clknet_1_0__leaf_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net862 (.A(clknet_0_net862),
    .X(clknet_1_1__leaf_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net638 (.A(net638),
    .X(clknet_0_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net638 (.A(clknet_0_net638),
    .X(clknet_1_0__leaf_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net638 (.A(clknet_0_net638),
    .X(clknet_1_1__leaf_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net637 (.A(net637),
    .X(clknet_0_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net637 (.A(clknet_0_net637),
    .X(clknet_1_0__leaf_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net637 (.A(clknet_0_net637),
    .X(clknet_1_1__leaf_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net390 (.A(net390),
    .X(clknet_0_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net390 (.A(clknet_0_net390),
    .X(clknet_1_0__leaf_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net390 (.A(clknet_0_net390),
    .X(clknet_1_1__leaf_net390));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net898 (.A(net898),
    .X(clknet_0_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net168 (.A(net168),
    .X(clknet_0_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_0__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_1__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net223 (.A(net223),
    .X(clknet_0_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_0__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_1__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net238 (.A(net238),
    .X(clknet_0_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net950 (.A(net950),
    .X(clknet_0_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net950 (.A(clknet_0_net950),
    .X(clknet_1_0__leaf_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net950 (.A(clknet_0_net950),
    .X(clknet_1_1__leaf_net950));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net970 (.A(net970),
    .X(clknet_0_net970));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net970 (.A(clknet_0_net970),
    .X(clknet_1_0__leaf_net970));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net970 (.A(clknet_0_net970),
    .X(clknet_1_1__leaf_net970));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net806 (.A(net806),
    .X(clknet_0_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net806 (.A(clknet_0_net806),
    .X(clknet_1_0__leaf_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net806 (.A(clknet_0_net806),
    .X(clknet_1_1__leaf_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net233 (.A(net233),
    .X(clknet_0_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net165 (.A(net165),
    .X(clknet_0_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net422 (.A(net422),
    .X(clknet_0_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_0__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_1__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net426 (.A(net426),
    .X(clknet_0_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net426 (.A(clknet_0_net426),
    .X(clknet_1_0__leaf_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net426 (.A(clknet_0_net426),
    .X(clknet_1_1__leaf_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net558 (.A(net558),
    .X(clknet_0_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_0__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net558 (.A(clknet_0_net558),
    .X(clknet_1_1__leaf_net558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net550 (.A(net550),
    .X(clknet_0_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_0__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_1__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net659 (.A(net659),
    .X(clknet_0_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net659 (.A(clknet_0_net659),
    .X(clknet_1_0__leaf_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net659 (.A(clknet_0_net659),
    .X(clknet_1_1__leaf_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net702 (.A(net702),
    .X(clknet_0_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_0__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_1__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net547 (.A(net547),
    .X(clknet_0_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net547 (.A(clknet_0_net547),
    .X(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net547 (.A(clknet_0_net547),
    .X(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net549 (.A(net549),
    .X(clknet_0_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_0__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_1__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net860 (.A(net860),
    .X(clknet_0_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net860 (.A(clknet_0_net860),
    .X(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net860 (.A(clknet_0_net860),
    .X(clknet_1_1__leaf_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net428 (.A(net428),
    .X(clknet_0_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net428 (.A(clknet_0_net428),
    .X(clknet_1_0__leaf_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net428 (.A(clknet_0_net428),
    .X(clknet_1_1__leaf_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net430 (.A(net430),
    .X(clknet_0_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net430 (.A(clknet_0_net430),
    .X(clknet_1_0__leaf_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net430 (.A(clknet_0_net430),
    .X(clknet_1_1__leaf_net430));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net295 (.A(net295),
    .X(clknet_0_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net313 (.A(net313),
    .X(clknet_0_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net313 (.A(clknet_0_net313),
    .X(clknet_1_0__leaf_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net313 (.A(clknet_0_net313),
    .X(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net171 (.A(net171),
    .X(clknet_0_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net171 (.A(clknet_0_net171),
    .X(clknet_1_0__leaf_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net171 (.A(clknet_0_net171),
    .X(clknet_1_1__leaf_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net585 (.A(net585),
    .X(clknet_0_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_0__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_1__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net587 (.A(net587),
    .X(clknet_0_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net587 (.A(clknet_0_net587),
    .X(clknet_1_0__leaf_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net587 (.A(clknet_0_net587),
    .X(clknet_1_1__leaf_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net576 (.A(net576),
    .X(clknet_0_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net576 (.A(clknet_0_net576),
    .X(clknet_1_0__leaf_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net576 (.A(clknet_0_net576),
    .X(clknet_1_1__leaf_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net589 (.A(net589),
    .X(clknet_0_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net589 (.A(clknet_0_net589),
    .X(clknet_1_0__leaf_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net589 (.A(clknet_0_net589),
    .X(clknet_1_1__leaf_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net167 (.A(net167),
    .X(clknet_0_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_0__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_1__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net435 (.A(net435),
    .X(clknet_0_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_0__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net561 (.A(net561),
    .X(clknet_0_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_0__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_1__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net557 (.A(net557),
    .X(clknet_0_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_0__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_1__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net170 (.A(net170),
    .X(clknet_0_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_0__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net170 (.A(clknet_0_net170),
    .X(clknet_1_1__leaf_net170));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net205 (.A(net205),
    .X(clknet_0_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_0__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net205 (.A(clknet_0_net205),
    .X(clknet_1_1__leaf_net205));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net331 (.A(net331),
    .X(clknet_0_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_0__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_1__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net823 (.A(net823),
    .X(clknet_0_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net463 (.A(net463),
    .X(clknet_0_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_0__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net463 (.A(clknet_0_net463),
    .X(clknet_1_1__leaf_net463));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net596 (.A(net596),
    .X(clknet_0_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_1__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net824 (.A(net824),
    .X(clknet_0_net824));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net824 (.A(clknet_0_net824),
    .X(clknet_1_0__leaf_net824));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net824 (.A(clknet_0_net824),
    .X(clknet_1_1__leaf_net824));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net369 (.A(net369),
    .X(clknet_0_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_0__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_1__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net358 (.A(net358),
    .X(clknet_0_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_0__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_1__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net966 (.A(net966),
    .X(clknet_0_net966));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net966 (.A(clknet_0_net966),
    .X(clknet_1_0__leaf_net966));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net966 (.A(clknet_0_net966),
    .X(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net958 (.A(net958),
    .X(clknet_0_net958));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net958 (.A(clknet_0_net958),
    .X(clknet_1_0__leaf_net958));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net958 (.A(clknet_0_net958),
    .X(clknet_1_1__leaf_net958));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net594 (.A(net594),
    .X(clknet_0_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net594 (.A(clknet_0_net594),
    .X(clknet_1_0__leaf_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net594 (.A(clknet_0_net594),
    .X(clknet_1_1__leaf_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net341 (.A(net341),
    .X(clknet_0_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_0__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net341 (.A(clknet_0_net341),
    .X(clknet_1_1__leaf_net341));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net207 (.A(net207),
    .X(clknet_0_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_0__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net211 (.A(net211),
    .X(clknet_0_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net211 (.A(clknet_0_net211),
    .X(clknet_1_0__leaf_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net211 (.A(clknet_0_net211),
    .X(clknet_1_1__leaf_net211));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net844 (.A(net844),
    .X(clknet_0_net844));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net844 (.A(clknet_0_net844),
    .X(clknet_1_0__leaf_net844));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net844 (.A(clknet_0_net844),
    .X(clknet_1_1__leaf_net844));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net198 (.A(net198),
    .X(clknet_0_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net202 (.A(net202),
    .X(clknet_0_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net213 (.A(net213),
    .X(clknet_0_net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net213 (.A(clknet_0_net213),
    .X(clknet_1_0__leaf_net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net213 (.A(clknet_0_net213),
    .X(clknet_1_1__leaf_net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net208 (.A(net208),
    .X(clknet_0_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_0__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net208 (.A(clknet_0_net208),
    .X(clknet_1_1__leaf_net208));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net897 (.A(net897),
    .X(clknet_0_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net398 (.A(net398),
    .X(clknet_0_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_0__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net398 (.A(clknet_0_net398),
    .X(clknet_1_1__leaf_net398));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net446 (.A(net446),
    .X(clknet_0_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_1__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net694 (.A(net694),
    .X(clknet_0_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net718 (.A(net718),
    .X(clknet_0_net718));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net718 (.A(clknet_0_net718),
    .X(clknet_1_0__leaf_net718));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net718 (.A(clknet_0_net718),
    .X(clknet_1_1__leaf_net718));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net593 (.A(net593),
    .X(clknet_0_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net593 (.A(clknet_0_net593),
    .X(clknet_1_0__leaf_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net593 (.A(clknet_0_net593),
    .X(clknet_1_1__leaf_net593));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net842 (.A(net842),
    .X(clknet_0_net842));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net842 (.A(clknet_0_net842),
    .X(clknet_1_0__leaf_net842));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net842 (.A(clknet_0_net842),
    .X(clknet_1_1__leaf_net842));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net586 (.A(net586),
    .X(clknet_0_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net586 (.A(clknet_0_net586),
    .X(clknet_1_0__leaf_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net586 (.A(clknet_0_net586),
    .X(clknet_1_1__leaf_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net405 (.A(net405),
    .X(clknet_0_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_0__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_1__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net395 (.A(net395),
    .X(clknet_0_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net395 (.A(clknet_0_net395),
    .X(clknet_1_0__leaf_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net395 (.A(clknet_0_net395),
    .X(clknet_1_1__leaf_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net416 (.A(net416),
    .X(clknet_0_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net416 (.A(clknet_0_net416),
    .X(clknet_1_0__leaf_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net416 (.A(clknet_0_net416),
    .X(clknet_1_1__leaf_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net431 (.A(net431),
    .X(clknet_0_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net431 (.A(clknet_0_net431),
    .X(clknet_1_0__leaf_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net431 (.A(clknet_0_net431),
    .X(clknet_1_1__leaf_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net425 (.A(net425),
    .X(clknet_0_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_0__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_1__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net432 (.A(net432),
    .X(clknet_0_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net432 (.A(clknet_0_net432),
    .X(clknet_1_0__leaf_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net432 (.A(clknet_0_net432),
    .X(clknet_1_1__leaf_net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net861 (.A(net861),
    .X(clknet_0_net861));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net861 (.A(clknet_0_net861),
    .X(clknet_1_0__leaf_net861));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net861 (.A(clknet_0_net861),
    .X(clknet_1_1__leaf_net861));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net946),
    .X(net154));
 sky130_fd_sc_hd__or2_1 clone2 (.A(net55),
    .B(net45),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(clknet_0_net602),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(clknet_0_net608),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net841),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net836),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net796),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net850),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net872),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net751),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net802),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net582),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net949),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net830),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net648),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net219),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net307),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net242),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net829),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net859),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net444),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net819),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(net38),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_1 wire2 (.A(net539),
    .X(net1032));
 sky130_fd_sc_hd__clkbuf_1 max_cap3 (.A(net661),
    .X(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_C1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A_N (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_Y (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A_N (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_S1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_D_N (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A_N (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_C_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_C_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_Y (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_S1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_Y (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_SCE (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_Y (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_Y (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_C1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_C1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_Y (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_RESET_B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B_N (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B_N (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A_N (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_Y (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_S0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_RESET_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_D1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_C1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_C (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_C (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B_N (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_C (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_Y (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_D_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_Y (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_S0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_D_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_S1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_D (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B_N (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SCD (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_C1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_S1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_C (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_S0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A_N (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_A3 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_Y (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_RESET_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A3 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_S1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_RESET_B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_SET_B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_SCE (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_D_N (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_Q_N (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_Q (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_Y (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_B_N (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_D_N (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_C_N (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S0 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_SCD (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_C_N (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_C_N (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_C (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_Y (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_RESET_B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_D (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_DE (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_C_N (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCE (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_SCE (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_Y (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_D_N (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_S1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_D_N (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_Y (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A3 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A3 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_C (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_Q_N (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_Q (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_SET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_D_N (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net198_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_Y (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_B_N (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_C_N (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_SCD (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_SCE (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_C (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_Y (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_C_N (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_Y (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_C1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_C_N (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_C_N (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_C (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B_N (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_RESET_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A3 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A3 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_X (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_S0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_D_N (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_C_N (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_SCE (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_D_N (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_S1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_Q_N (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_S0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_C_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_C_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_Q (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A3 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_C_N (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A_N (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_Y (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S0 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_SCE (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_C_N (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_D1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_D_N (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_Y (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_C (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_SET_B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_Y (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B_N (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_C_N (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_C1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_C (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_C_N (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_C_N (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_SCE (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_C_N (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_C (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_Y (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_X (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SCD (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_SCD (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_Y (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net295_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_Y (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_C1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_D (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A0 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_C (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_S0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_C_N (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_SCD (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_D_N (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_C1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_C_N (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A3 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B_N (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_B (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_Y (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A3 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_C (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold17_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_D (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_Y (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_S0 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A0 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_SCD (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_SCD (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_Y (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_X (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_X (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_Y (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_D_N (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A0 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_C_N (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_Y (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_Q (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c60_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_D (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Y (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A3 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_S0 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_C1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_RESET_B (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S0 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Y (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_S0 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_SCD (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SCE (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_D1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SCD (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A_N (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SCE (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_Y (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_D (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_D (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_Y (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_SCD (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_B_N (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_D (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A1 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_Q (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A_N (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_S0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A_N (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap76_A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_D (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_C_N (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_C (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_B (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_Y (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_B1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_C1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_RESET_B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_SCD (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_Y (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_Y (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_D_N (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_Q_N (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCD (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_RESET_B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_Q (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_Q (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A_N (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A0 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_D (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_B (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_D (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_Y (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A3 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_C_N (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A1 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_Y (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A0 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_X (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net529_A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_X (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A3 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A0 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B_N (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_Y (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_S1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A0 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_SET_B (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_C_N (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_X (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_B1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_C_N (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A0 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_X (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_Y (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_D (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_SCD (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_S0 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_SCE (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_RESET_B (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_B1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_D1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCE (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A_N (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_B (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_X (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_X (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A_N (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_Y (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_B1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_D (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A3 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_X (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_C1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_Q_N (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_C (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_Q (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A3 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_SCE (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_D1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_B1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_Q (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_X (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_C_N (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_B (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_Q_N (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A0 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_SCD (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_Q (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_X (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_D1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_Y (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A3 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_C1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_X (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold15_A (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_D1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_B1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_Y (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_S0 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_SCE (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_B1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_X (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_X (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_RESET_B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_C_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_Q (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_S1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_Q_N (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_SCD (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_Q (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_SET_B (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_SCE (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_D_N (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_B (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_SCE (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_Y (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_Q (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_D1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B_N (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_B (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_D1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B_N (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_B (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_C_N (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_RESET_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A_N (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_D1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_s844_Q (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_S1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_SCE (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_SET_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_S1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_D_N (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_s849_Q (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_D1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_Q (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_D1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_D1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_D1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_B (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_Q (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_S1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_S1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_C_N (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_C (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_C (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_C_N (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_Q (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_D1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_S0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A_N (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_SET_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_S0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_B_N (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B_N (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_Q (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SET_B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_D1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SCE (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_D1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_C_N (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_C (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_Q (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net861_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_GCLK (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_Q (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net898_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_GCLK (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_RESET_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_A_N (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_Y (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_C1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_Q (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_Q (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_RESET_B (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B_N (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SCE (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_SET_B (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_B (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_A_N (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B_N (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_B (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B_N (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_C (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A_N (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_SCE (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_B (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_C1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C_N (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B_N (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_B (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_D1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_C (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_B (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_B (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A2 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_C (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A_N (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_C (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_D (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B_N (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_D_N (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A_N (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_C1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_C (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_RESET_B (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_X (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_C1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_B1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_RESET_B (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_Y (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold13_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_B1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_SCD (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_B1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_B1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_S1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_SCD (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_D1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_SCE (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCD (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_SCE (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_SET_B (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_C1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_D (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_SCE (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_B1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_SCE (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_SCD (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_SCE (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_D1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_C_N (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_D1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_B (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_DE (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_C_N (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap62_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_SET_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_C_N (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCE (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_C (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_C1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_SCD (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_C (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_B (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_C (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_C1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_C (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_B1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_D1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap66_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_C (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A_N (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_C_N (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_C1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_C (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_C (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_C (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_C (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B_N (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_D_N (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_D1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B_N (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_D1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_C (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A2 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_D1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_C (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_C1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_C_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_C1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_D1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_C_N (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_B1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_SCE (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_D_N (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap76_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B_N (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_SCD (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_B1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_C_N (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_B_N (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_C_N (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_SCE (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_SET_B (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCE (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_C (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_C (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_C1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_D_N (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s843_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_SLEEP_B (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s845_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s846_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s842_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s850_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s844_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s847_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s848_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s851_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_B (.DIODE(clknet_1_0__leaf_net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(clknet_1_0__leaf_net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A2 (.DIODE(clknet_1_0__leaf_net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net634_X (.DIODE(clknet_1_0__leaf_net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S1 (.DIODE(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_C1 (.DIODE(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net951_X (.DIODE(clknet_1_1__leaf_net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net529_A (.DIODE(clknet_0_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net529_A (.DIODE(clknet_0_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net529_X (.DIODE(clknet_0_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A3 (.DIODE(clknet_1_0__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(clknet_1_0__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_D_N (.DIODE(clknet_1_0__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A1 (.DIODE(clknet_1_0__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net529_X (.DIODE(clknet_1_0__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_RESET_B (.DIODE(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net529_X (.DIODE(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_1_A (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_net999_2_A (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_5_A (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_6_A (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_7_A (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net898_X (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B (.DIODE(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_D_N (.DIODE(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_SCE (.DIODE(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_D_N (.DIODE(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S1 (.DIODE(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net547_X (.DIODE(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net547_X (.DIODE(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_D1 (.DIODE(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_D_N (.DIODE(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A1 (.DIODE(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A2 (.DIODE(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_S0 (.DIODE(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net295_X (.DIODE(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_S1 (.DIODE(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A3 (.DIODE(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A0 (.DIODE(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net295_X (.DIODE(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S1 (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S1 (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_SCE (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net823_X (.DIODE(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_S0 (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_SET_B (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_SET_B (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net823_X (.DIODE(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(clknet_1_0__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SET_B (.DIODE(clknet_1_0__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_D1 (.DIODE(clknet_1_0__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_B1 (.DIODE(clknet_1_0__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(clknet_1_0__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net958_X (.DIODE(clknet_1_0__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_S1 (.DIODE(clknet_1_1__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_D1 (.DIODE(clknet_1_1__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_S1 (.DIODE(clknet_1_1__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(clknet_1_1__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net958_X (.DIODE(clknet_1_1__leaf_net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_C (.DIODE(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_SCE (.DIODE(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_RESET_B (.DIODE(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net198_X (.DIODE(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net198_X (.DIODE(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_D_N (.DIODE(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_SCE (.DIODE(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net446_X (.DIODE(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_X (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold13_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net125));
 sky130_fd_sc_hd__or2_1 clone1 (.A(net45),
    .B(net55),
    .X(net1034));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
