module netlist_2 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire clknet_0_clk;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net678;
 wire clknet_1_0__leaf_net678;
 wire clknet_1_1__leaf_net678;
 wire clknet_0_net596;
 wire clknet_1_0__leaf_net596;
 wire clknet_1_1__leaf_net596;
 wire clknet_0_net594;
 wire clknet_1_0__leaf_net594;
 wire clknet_1_1__leaf_net594;
 wire clknet_0_net496;
 wire clknet_1_0__leaf_net496;
 wire clknet_1_1__leaf_net496;
 wire clknet_0_net505;
 wire clknet_1_0__leaf_net505;
 wire clknet_1_1__leaf_net505;
 wire clknet_0_net517;
 wire clknet_1_0__leaf_net517;
 wire clknet_1_1__leaf_net517;
 wire clknet_0_net499;
 wire clknet_1_0__leaf_net499;
 wire clknet_1_1__leaf_net499;
 wire clknet_0_net676;
 wire clknet_1_0__leaf_net676;
 wire clknet_1_1__leaf_net676;
 wire clknet_0_net677;
 wire clknet_1_0__leaf_net677;
 wire clknet_1_1__leaf_net677;
 wire clknet_0_net526;
 wire clknet_1_0__leaf_net526;
 wire clknet_1_1__leaf_net526;
 wire clknet_0_net521;
 wire clknet_1_0__leaf_net521;
 wire clknet_1_1__leaf_net521;
 wire clknet_0_net497;
 wire clknet_1_0__leaf_net497;
 wire clknet_1_1__leaf_net497;
 wire clknet_0_net504;
 wire clknet_1_0__leaf_net504;
 wire clknet_1_1__leaf_net504;
 wire clknet_0_net513;
 wire clknet_1_0__leaf_net513;
 wire clknet_1_1__leaf_net513;
 wire clknet_0_net657;
 wire clknet_1_0__leaf_net657;
 wire clknet_1_1__leaf_net657;
 wire clknet_0_net656;
 wire clknet_1_0__leaf_net656;
 wire clknet_1_1__leaf_net656;
 wire clknet_0_net423;
 wire clknet_1_0__leaf_net423;
 wire clknet_1_1__leaf_net423;
 wire clknet_0_net655;
 wire clknet_1_0__leaf_net655;
 wire clknet_1_1__leaf_net655;
 wire clknet_0_net418;
 wire clknet_1_0__leaf_net418;
 wire clknet_1_1__leaf_net418;
 wire clknet_0_net637;
 wire clknet_1_0__leaf_net637;
 wire clknet_1_1__leaf_net637;
 wire clknet_0_net404;
 wire clknet_1_0__leaf_net404;
 wire clknet_1_1__leaf_net404;
 wire clknet_0_net393;
 wire clknet_1_0__leaf_net393;
 wire clknet_1_1__leaf_net393;
 wire clknet_0_net377;
 wire clknet_1_0__leaf_net377;
 wire clknet_1_1__leaf_net377;
 wire clknet_0_net378;
 wire clknet_1_0__leaf_net378;
 wire clknet_1_1__leaf_net378;
 wire clknet_0_net636;
 wire clknet_1_0__leaf_net636;
 wire clknet_1_1__leaf_net636;
 wire clknet_0_net635;
 wire clknet_1_0__leaf_net635;
 wire clknet_1_1__leaf_net635;
 wire clknet_0_net803;
 wire clknet_1_0__leaf_net803;
 wire clknet_1_1__leaf_net803;
 wire clknet_0_net617;
 wire clknet_1_0__leaf_net617;
 wire clknet_1_1__leaf_net617;
 wire clknet_0_net807;
 wire clknet_1_0__leaf_net807;
 wire clknet_1_1__leaf_net807;
 wire clknet_0_net798;
 wire clknet_1_0__leaf_net798;
 wire clknet_1_1__leaf_net798;
 wire clknet_0_net616;
 wire clknet_1_0__leaf_net616;
 wire clknet_1_1__leaf_net616;
 wire clknet_0_net834;
 wire clknet_1_0__leaf_net834;
 wire clknet_1_1__leaf_net834;
 wire clknet_0_net822;
 wire clknet_1_0__leaf_net822;
 wire clknet_1_1__leaf_net822;
 wire clknet_0_net200;
 wire clknet_1_0__leaf_net200;
 wire clknet_1_1__leaf_net200;
 wire clknet_0_net840;
 wire clknet_1_0__leaf_net840;
 wire clknet_1_1__leaf_net840;
 wire clknet_0_net309;
 wire clknet_1_0__leaf_net309;
 wire clknet_1_1__leaf_net309;
 wire clknet_0_net303;
 wire clknet_1_0__leaf_net303;
 wire clknet_1_1__leaf_net303;
 wire clknet_0_net189;
 wire clknet_1_0__leaf_net189;
 wire clknet_1_1__leaf_net189;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net483;
 wire clknet_1_0__leaf_net483;
 wire clknet_1_1__leaf_net483;
 wire clknet_0_net472;
 wire clknet_1_0__leaf_net472;
 wire clknet_1_1__leaf_net472;
 wire clknet_0_net355;
 wire clknet_1_0__leaf_net355;
 wire clknet_1_1__leaf_net355;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire net442;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;

 sky130_fd_sc_hd__a41oi_2 c100 (.A1(net779),
    .A2(net886),
    .A3(net889),
    .A4(net780),
    .B1(net771),
    .Y(net0));
 sky130_fd_sc_hd__mux4_2 c101 (.A0(net771),
    .A1(net777),
    .A2(net0),
    .A3(net776),
    .S0(net889),
    .S1(net886),
    .X(net1));
 sky130_fd_sc_hd__a41oi_4 c102 (.A1(net774),
    .A2(net1),
    .A3(net764),
    .A4(net766),
    .B1(net727),
    .Y(net2));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net722),
    .A1(net711),
    .A2(net2),
    .A3(net775),
    .S0(net781),
    .S1(net892),
    .X(net3));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net711),
    .A1(net2),
    .A2(net773),
    .A3(net722),
    .S0(net889),
    .S1(net777),
    .X(net837));
 sky130_fd_sc_hd__mux4_2 c105 (.A0(net1),
    .A1(net781),
    .A2(net779),
    .A3(net771),
    .S0(net889),
    .S1(net3),
    .X(net847));
 sky130_fd_sc_hd__a41o_1 c106 (.A1(net2),
    .A2(net777),
    .A3(net764),
    .A4(net847),
    .B1(net886),
    .X(net4));
 sky130_fd_sc_hd__mux4_2 c107 (.A0(net837),
    .A1(net3),
    .A2(net705),
    .A3(net1),
    .S0(net773),
    .S1(net847),
    .X(net5));
 sky130_fd_sc_hd__mux4_2 c108 (.A0(net5),
    .A1(net837),
    .A2(net756),
    .A3(net889),
    .S0(net3),
    .S1(net847),
    .X(net851));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net4),
    .A1(net3),
    .A2(net773),
    .A3(net718),
    .S0(net774),
    .S1(net837),
    .X(net852));
 sky130_fd_sc_hd__mux4_2 c122 (.A0(net703),
    .A1(net782),
    .A2(net747),
    .A3(net748),
    .S0(net5),
    .S1(net779),
    .X(net831));
 sky130_fd_sc_hd__mux4_2 c123 (.A0(net5),
    .A1(net831),
    .A2(net837),
    .A3(net847),
    .S0(net851),
    .S1(net715),
    .X(net842));
 sky130_fd_sc_hd__a41o_1 c124 (.A1(net842),
    .A2(net2),
    .A3(net851),
    .A4(net715),
    .B1(net779),
    .X(net6));
 sky130_fd_sc_hd__mux4_2 c125 (.A0(net748),
    .A1(net6),
    .A2(net744),
    .A3(net852),
    .S0(net837),
    .S1(net725),
    .X(net849));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net6),
    .A1(net849),
    .A2(net718),
    .A3(net847),
    .S0(net831),
    .S1(net842),
    .X(net854));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net6),
    .A1(net849),
    .A2(net842),
    .A3(net851),
    .S0(net887),
    .S1(net854),
    .X(net855));
 sky130_fd_sc_hd__mux4_2 c128 (.A0(net855),
    .A1(net831),
    .A2(net842),
    .A3(net6),
    .S0(net778),
    .S1(net849),
    .X(net846));
 sky130_fd_sc_hd__mux4_2 c129 (.A0(net854),
    .A1(net1),
    .A2(net846),
    .A3(net6),
    .S0(net837),
    .S1(net756),
    .X(net850));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net738),
    .A1(net846),
    .A2(net855),
    .A3(net849),
    .S0(net850),
    .S1(net6),
    .X(net853));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net715),
    .A1(net853),
    .A2(net855),
    .A3(net850),
    .S0(net849),
    .S1(net6),
    .X(net7));
 sky130_fd_sc_hd__a21boi_4 c132 (.A1(net707),
    .A2(net761),
    .B1_N(net890),
    .Y(net8));
 sky130_fd_sc_hd__xnor2_4 c133 (.A(net729),
    .B(net8),
    .Y(net9));
 sky130_fd_sc_hd__xor2_4 c134 (.A(net688),
    .B(net707),
    .X(net10));
 sky130_fd_sc_hd__xor2_4 c135 (.A(net750),
    .B(net707),
    .X(net11));
 sky130_fd_sc_hd__a21oi_4 c136 (.A1(net691),
    .A2(net884),
    .B1(net688),
    .Y(net12));
 sky130_fd_sc_hd__o21ba_2 c137 (.A1(net687),
    .A2(net690),
    .B1_N(net890),
    .X(net13));
 sky130_fd_sc_hd__o21ai_4 c138 (.A1(net12),
    .A2(net13),
    .B1(net890),
    .Y(net14));
 sky130_fd_sc_hd__xor2_4 c139 (.A(net698),
    .B(net750),
    .X(net15));
 sky130_fd_sc_hd__a41oi_4 c140 (.A1(net693),
    .A2(net696),
    .A3(net11),
    .A4(net15),
    .B1(net884),
    .Y(net16));
 sky130_fd_sc_hd__a21oi_4 c141 (.A1(net13),
    .A2(net690),
    .B1(net16),
    .Y(net17));
 sky130_fd_sc_hd__a41o_2 c142 (.A1(net686),
    .A2(net14),
    .A3(net906),
    .A4(net16),
    .B1(net9),
    .X(net18));
 sky130_fd_sc_hd__o21ai_4 c143 (.A1(net739),
    .A2(net9),
    .B1(net15),
    .Y(net19));
 sky130_fd_sc_hd__mux2_4 c144 (.A0(net16),
    .A1(net890),
    .S(net17),
    .X(net20));
 sky130_fd_sc_hd__a21o_1 c145 (.A1(net9),
    .A2(net884),
    .B1(net18),
    .X(net21));
 sky130_fd_sc_hd__a21oi_1 c146 (.A1(net11),
    .A2(net21),
    .B1(net14),
    .Y(net22));
 sky130_fd_sc_hd__a21bo_4 c147 (.A1(net20),
    .A2(net16),
    .B1_N(net884),
    .X(net23));
 sky130_fd_sc_hd__o21ba_2 c148 (.A1(net21),
    .A2(net18),
    .B1_N(net688),
    .X(net24));
 sky130_fd_sc_hd__a41oi_4 c149 (.A1(net14),
    .A2(net24),
    .A3(net750),
    .A4(net21),
    .B1(net697),
    .Y(net25));
 sky130_fd_sc_hd__mux2_2 c150 (.A0(net697),
    .A1(net25),
    .S(net693),
    .X(net26));
 sky130_fd_sc_hd__mux4_1 c151 (.A0(net18),
    .A1(net23),
    .A2(net26),
    .A3(net15),
    .S0(net22),
    .S1(net690),
    .X(net27));
 sky130_fd_sc_hd__o21ai_2 c152 (.A1(net27),
    .A2(net25),
    .B1(net23),
    .Y(net28));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net15),
    .A1(net28),
    .A2(net20),
    .A3(net13),
    .S0(net25),
    .S1(net23),
    .X(net841));
 sky130_fd_sc_hd__a21oi_4 c154 (.A1(net694),
    .A2(net871),
    .B1(net710),
    .Y(net29));
 sky130_fd_sc_hd__o21ai_4 c155 (.A1(net719),
    .A2(net709),
    .B1(net702),
    .Y(net30));
 sky130_fd_sc_hd__mux2_4 c156 (.A0(net702),
    .A1(net709),
    .S(net714),
    .X(net31));
 sky130_fd_sc_hd__a31o_2 c157 (.A1(net721),
    .A2(net31),
    .A3(net701),
    .B1(net99),
    .X(net32));
 sky130_fd_sc_hd__o21ba_1 c158 (.A1(net27),
    .A2(net702),
    .B1_N(net714),
    .X(net33));
 sky130_fd_sc_hd__a21oi_2 c159 (.A1(net30),
    .A2(net717),
    .B1(net32),
    .Y(net34));
 sky130_fd_sc_hd__mux2_2 c160 (.A0(net26),
    .A1(net33),
    .S(net717),
    .X(net35));
 sky130_fd_sc_hd__a21oi_4 c161 (.A1(net13),
    .A2(net692),
    .B1(net702),
    .Y(net36));
 sky130_fd_sc_hd__a31oi_4 c162 (.A1(net717),
    .A2(net701),
    .A3(net714),
    .B1(net26),
    .Y(net843));
 sky130_fd_sc_hd__a21o_1 c163 (.A1(net843),
    .A2(net32),
    .B1(net24),
    .X(net37));
 sky130_fd_sc_hd__o21a_4 c164 (.A1(net36),
    .A2(net713),
    .B1(net31),
    .X(net825));
 sky130_fd_sc_hd__a31o_1 c165 (.A1(net35),
    .A2(net34),
    .A3(net825),
    .B1(net843),
    .X(net38));
 sky130_fd_sc_hd__a31oi_2 c166 (.A1(net720),
    .A2(net31),
    .A3(net38),
    .B1(net843),
    .Y(net39));
 sky130_fd_sc_hd__a41o_1 c167 (.A1(net22),
    .A2(net31),
    .A3(net38),
    .A4(net843),
    .B1(net30),
    .X(net40));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net39),
    .A1(net14),
    .A2(net32),
    .A3(net35),
    .S0(net13),
    .S1(net703),
    .X(net41));
 sky130_fd_sc_hd__a31o_1 c169 (.A1(net38),
    .A2(net33),
    .A3(net30),
    .B1(net861),
    .X(net42));
 sky130_fd_sc_hd__mux4_1 c170 (.A0(net36),
    .A1(net843),
    .A2(net42),
    .A3(net40),
    .S0(net30),
    .S1(net861),
    .X(net43));
 sky130_fd_sc_hd__a21boi_2 c171 (.A1(net710),
    .A2(net692),
    .B1_N(net566),
    .Y(net44));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net42),
    .A1(net712),
    .A2(net44),
    .A3(net714),
    .S0(net861),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net33),
    .A1(net40),
    .A2(net825),
    .A3(net37),
    .S0(net26),
    .S1(net567),
    .X(net46));
 sky130_fd_sc_hd__a31oi_1 c174 (.A1(net44),
    .A2(net39),
    .A3(net861),
    .B1(net567),
    .Y(net47));
 sky130_fd_sc_hd__mux2_2 c175 (.A0(net37),
    .A1(net46),
    .S(net704),
    .X(net795));
 sky130_fd_sc_hd__a21boi_4 c176 (.A1(net726),
    .A2(net30),
    .B1_N(net703),
    .Y(net48));
 sky130_fd_sc_hd__o21ai_2 c177 (.A1(net32),
    .A2(net734),
    .B1(net725),
    .Y(net49));
 sky130_fd_sc_hd__a31o_1 c178 (.A1(net728),
    .A2(net48),
    .A3(net734),
    .B1(net705),
    .X(net50));
 sky130_fd_sc_hd__a41oi_4 c179 (.A1(net825),
    .A2(net724),
    .A3(net48),
    .A4(net706),
    .B1(net692),
    .Y(net814));
 sky130_fd_sc_hd__a41oi_2 c180 (.A1(net731),
    .A2(net50),
    .A3(net724),
    .A4(net745),
    .B1(net895),
    .Y(net51));
 sky130_fd_sc_hd__a31o_4 c181 (.A1(net23),
    .A2(net737),
    .A3(net706),
    .B1(net895),
    .X(net52));
 sky130_fd_sc_hd__a41o_2 c182 (.A1(net699),
    .A2(net692),
    .A3(net34),
    .A4(net874),
    .B1(net49),
    .X(net53));
 sky130_fd_sc_hd__a31oi_2 c183 (.A1(net50),
    .A2(net723),
    .A3(net32),
    .B1(net872),
    .Y(net54));
 sky130_fd_sc_hd__a21bo_2 c184 (.A1(net740),
    .A2(net880),
    .B1_N(net51),
    .X(net55));
 sky130_fd_sc_hd__a41oi_4 c185 (.A1(net52),
    .A2(net712),
    .A3(net23),
    .A4(net731),
    .B1(net890),
    .Y(net56));
 sky130_fd_sc_hd__a41o_1 c186 (.A1(net870),
    .A2(net50),
    .A3(net49),
    .A4(net736),
    .B1(net872),
    .X(net57));
 sky130_fd_sc_hd__a41oi_4 c187 (.A1(net35),
    .A2(net700),
    .A3(net52),
    .A4(net872),
    .B1(net903),
    .Y(net58));
 sky130_fd_sc_hd__mux4_2 c188 (.A0(net734),
    .A1(net57),
    .A2(net723),
    .A3(net870),
    .S0(net874),
    .S1(net872),
    .X(net59));
 sky130_fd_sc_hd__a41o_1 c189 (.A1(net723),
    .A2(net874),
    .A3(net903),
    .A4(net872),
    .B1(net58),
    .X(net60));
 sky130_fd_sc_hd__mux4_1 c190 (.A0(net54),
    .A1(net58),
    .A2(net55),
    .A3(net59),
    .S0(net734),
    .S1(net60),
    .X(net61));
 sky130_fd_sc_hd__mux4_1 c191 (.A0(net872),
    .A1(net49),
    .A2(net54),
    .A3(net60),
    .S0(net48),
    .S1(net950),
    .X(net62));
 sky130_fd_sc_hd__a41oi_2 c192 (.A1(net24),
    .A2(net874),
    .A3(net62),
    .A4(net35),
    .B1(net728),
    .Y(net63));
 sky130_fd_sc_hd__mux4_1 c193 (.A0(net62),
    .A1(net55),
    .A2(net63),
    .A3(net700),
    .S0(net901),
    .S1(net723),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net57),
    .A1(net884),
    .A2(net737),
    .A3(net706),
    .S0(net734),
    .S1(net951),
    .X(net65));
 sky130_fd_sc_hd__mux4_4 c195 (.A0(net65),
    .A1(net858),
    .A2(net60),
    .A3(net725),
    .S0(net872),
    .S1(net592),
    .X(net66));
 sky130_fd_sc_hd__a41oi_1 c196 (.A1(net60),
    .A2(net54),
    .A3(net65),
    .A4(net858),
    .B1(net58),
    .Y(net67));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net61),
    .A1(net883),
    .A2(net734),
    .A3(net58),
    .S0(net858),
    .S1(net835),
    .X(net68));
 sky130_fd_sc_hd__o21ai_1 c198 (.A1(net741),
    .A2(net903),
    .B1(net759),
    .Y(net69));
 sky130_fd_sc_hd__mux2_4 c199 (.A0(net59),
    .A1(net889),
    .S(net887),
    .X(net839));
 sky130_fd_sc_hd__a31oi_1 c200 (.A1(net741),
    .A2(net701),
    .A3(net892),
    .B1(net835),
    .Y(net70));
 sky130_fd_sc_hd__a21o_4 c201 (.A1(net751),
    .A2(net839),
    .B1(net889),
    .X(net804));
 sky130_fd_sc_hd__o21bai_4 c202 (.A1(net749),
    .A2(net716),
    .B1_N(net591),
    .Y(net71));
 sky130_fd_sc_hd__o21ba_1 c203 (.A1(net753),
    .A2(net752),
    .B1_N(net59),
    .X(net72));
 sky130_fd_sc_hd__a41o_2 c204 (.A1(net70),
    .A2(net726),
    .A3(net895),
    .A4(net71),
    .B1(net72),
    .X(net786));
 sky130_fd_sc_hd__o21ba_2 c205 (.A1(net759),
    .A2(net71),
    .B1_N(net767),
    .X(net73));
 sky130_fd_sc_hd__a41o_4 c206 (.A1(net839),
    .A2(net701),
    .A3(net742),
    .A4(net754),
    .B1(net73),
    .X(net74));
 sky130_fd_sc_hd__a21bo_4 c207 (.A1(net74),
    .A2(net34),
    .B1_N(net72),
    .X(net844));
 sky130_fd_sc_hd__xor2_1 c208 (.A(net72),
    .B(net755),
    .X(net75));
 sky130_fd_sc_hd__mux4_2 c209 (.A0(net71),
    .A1(net839),
    .A2(net843),
    .A3(net73),
    .S0(net759),
    .S1(net874),
    .X(net76));
 sky130_fd_sc_hd__mux2_4 c210 (.A0(net767),
    .A1(net887),
    .S(net835),
    .X(net77));
 sky130_fd_sc_hd__a21boi_1 c211 (.A1(net844),
    .A2(net59),
    .B1_N(net872),
    .Y(net78));
 sky130_fd_sc_hd__a41oi_1 c212 (.A1(net69),
    .A2(net769),
    .A3(net76),
    .A4(net843),
    .B1(net751),
    .Y(net79));
 sky130_fd_sc_hd__o21ba_1 c213 (.A1(net757),
    .A2(net839),
    .B1_N(net76),
    .X(net80));
 sky130_fd_sc_hd__mux4_2 c214 (.A0(net75),
    .A1(net71),
    .A2(net74),
    .A3(net844),
    .S0(net77),
    .S1(net887),
    .X(net81));
 sky130_fd_sc_hd__mux4_2 c215 (.A0(net79),
    .A1(net10),
    .A2(net804),
    .A3(net81),
    .S0(net889),
    .S1(net73),
    .X(net827));
 sky130_fd_sc_hd__mux4_2 c216 (.A0(net742),
    .A1(net81),
    .A2(net78),
    .A3(net741),
    .S0(net71),
    .S1(net591),
    .X(net82));
 sky130_fd_sc_hd__a41o_1 c217 (.A1(net80),
    .A2(net73),
    .A3(net889),
    .A4(net752),
    .B1(net82),
    .X(net83));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net82),
    .A1(net81),
    .A2(net827),
    .A3(net76),
    .S0(net34),
    .S1(net592),
    .X(net84));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net83),
    .A1(net61),
    .A2(net81),
    .A3(net887),
    .S0(net827),
    .S1(net566),
    .X(net85));
 sky130_fd_sc_hd__a21oi_2 c220 (.A1(net718),
    .A2(net781),
    .B1(net743),
    .Y(net86));
 sky130_fd_sc_hd__o21ai_2 c221 (.A1(net773),
    .A2(net758),
    .B1(net74),
    .Y(net826));
 sky130_fd_sc_hd__o21ai_4 c222 (.A1(net889),
    .A2(net779),
    .B1(net778),
    .Y(net813));
 sky130_fd_sc_hd__mux4_2 c223 (.A0(net781),
    .A1(net82),
    .A2(net844),
    .A3(net874),
    .S0(net747),
    .S1(net883),
    .X(net87));
 sky130_fd_sc_hd__a21oi_2 c224 (.A1(net813),
    .A2(net743),
    .B1(net592),
    .Y(net88));
 sky130_fd_sc_hd__o21bai_4 c225 (.A1(net955),
    .A2(net902),
    .B1_N(net709),
    .Y(net823));
 sky130_fd_sc_hd__inv_6 c226 (.A(net574),
    .Y(net89));
 sky130_fd_sc_hd__a31oi_1 c227 (.A1(net775),
    .A2(net823),
    .A3(net827),
    .B1(net917),
    .Y(net90));
 sky130_fd_sc_hd__a21o_2 c228 (.A1(net813),
    .A2(net88),
    .B1(net887),
    .X(net91));
 sky130_fd_sc_hd__mux4_2 c229 (.A0(net730),
    .A1(net89),
    .A2(net88),
    .A3(net777),
    .S0(net763),
    .S1(net574),
    .X(net838));
 sky130_fd_sc_hd__a21bo_4 c230 (.A1(net727),
    .A2(net91),
    .B1_N(net89),
    .X(net92));
 sky130_fd_sc_hd__a41o_1 c231 (.A1(net780),
    .A2(net774),
    .A3(net89),
    .A4(net92),
    .B1(net827),
    .X(net93));
 sky130_fd_sc_hd__a41o_4 c232 (.A1(net0),
    .A2(net89),
    .A3(net774),
    .A4(net88),
    .B1(net838),
    .X(net94));
 sky130_fd_sc_hd__a41oi_4 c233 (.A1(net776),
    .A2(net86),
    .A3(net94),
    .A4(net813),
    .B1(net92),
    .Y(net95));
 sky130_fd_sc_hd__a31oi_2 c234 (.A1(net86),
    .A2(net89),
    .A3(net782),
    .B1(net779),
    .Y(net96));
 sky130_fd_sc_hd__a41o_1 c235 (.A1(net737),
    .A2(net92),
    .A3(net87),
    .A4(net838),
    .B1(net96),
    .X(net97));
 sky130_fd_sc_hd__a31o_4 c236 (.A1(net96),
    .A2(net92),
    .A3(net592),
    .B1(net845),
    .X(net817));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net96),
    .A1(net856),
    .A2(net74),
    .A3(net838),
    .S0(net89),
    .S1(net845),
    .X(net98));
 sky130_fd_sc_hd__mux4_2 c238 (.A0(net89),
    .A1(net87),
    .A2(net98),
    .A3(net866),
    .S0(net908),
    .X(net845));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net98),
    .A1(net826),
    .A2(net86),
    .A3(net94),
    .S0(net574),
    .S1(net845),
    .X(net100));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net100),
    .A1(net838),
    .A2(net856),
    .A3(net777),
    .S0(net89),
    .S1(net900),
    .X(net101));
 sky130_fd_sc_hd__mux4_2 c241 (.A0(net101),
    .A1(net98),
    .A2(net96),
    .A3(net763),
    .S0(net908),
    .S1(net100),
    .X(net818));
 sky130_fd_sc_hd__o21bai_4 c264 (.A1(net18),
    .A2(net99),
    .B1_N(net906),
    .Y(net102));
 sky130_fd_sc_hd__a21o_4 c265 (.A1(net102),
    .A2(net772),
    .B1(net906),
    .X(net103));
 sky130_fd_sc_hd__a21oi_4 c266 (.A1(net9),
    .A2(net102),
    .B1(net692),
    .Y(net104));
 sky130_fd_sc_hd__a21oi_4 c267 (.A1(net14),
    .A2(net20),
    .B1(net12),
    .Y(net105));
 sky130_fd_sc_hd__a21o_4 c268 (.A1(net102),
    .A2(net17),
    .B1(net28),
    .X(net106));
 sky130_fd_sc_hd__a21bo_2 c269 (.A1(net102),
    .A2(net18),
    .B1_N(net104),
    .X(net107));
 sky130_fd_sc_hd__mux2_4 c270 (.A0(net750),
    .A1(net105),
    .S(net685),
    .X(net108));
 sky130_fd_sc_hd__o21bai_4 c271 (.A1(net107),
    .A2(net105),
    .B1_N(net750),
    .Y(net109));
 sky130_fd_sc_hd__a21boi_4 c272 (.A1(net104),
    .A2(net103),
    .B1_N(net106),
    .Y(net110));
 sky130_fd_sc_hd__a31oi_4 c273 (.A1(net107),
    .A2(net105),
    .A3(net102),
    .B1(net9),
    .Y(net111));
 sky130_fd_sc_hd__o21ai_4 c274 (.A1(net111),
    .A2(net104),
    .B1(net906),
    .Y(net788));
 sky130_fd_sc_hd__xnor2_4 c275 (.A(net103),
    .B(net99),
    .Y(net112));
 sky130_fd_sc_hd__a21boi_4 c276 (.A1(net104),
    .A2(net110),
    .B1_N(net28),
    .Y(net113));
 sky130_fd_sc_hd__o21ba_4 c277 (.A1(net105),
    .A2(net109),
    .B1_N(net113),
    .X(net114));
 sky130_fd_sc_hd__mux4_2 c278 (.A0(net112),
    .A1(net106),
    .A2(net685),
    .A3(net103),
    .S0(net948),
    .S1(net18),
    .X(net115));
 sky130_fd_sc_hd__a41oi_4 c279 (.A1(net107),
    .A2(net113),
    .A3(net11),
    .A4(net104),
    .B1(net111),
    .Y(net116));
 sky130_fd_sc_hd__mux2_4 c280 (.A0(net110),
    .A1(net115),
    .S(net108),
    .X(net117));
 sky130_fd_sc_hd__mux4_2 c281 (.A0(net111),
    .A1(net115),
    .A2(net692),
    .A3(net108),
    .S0(net867),
    .S1(net113),
    .X(net794));
 sky130_fd_sc_hd__o21bai_4 c282 (.A1(net772),
    .A2(net11),
    .B1_N(net114),
    .Y(net832));
 sky130_fd_sc_hd__a31oi_1 c283 (.A1(net114),
    .A2(net832),
    .A3(net772),
    .B1(net112),
    .Y(net118));
 sky130_fd_sc_hd__a41o_1 c284 (.A1(net788),
    .A2(net112),
    .A3(net832),
    .A4(net106),
    .X(net119));
 sky130_fd_sc_hd__a21o_4 c285 (.A1(net117),
    .A2(net110),
    .B1(net116),
    .X(net120));
 sky130_fd_sc_hd__a21o_1 c286 (.A1(net102),
    .A2(net14),
    .B1(net701),
    .X(net121));
 sky130_fd_sc_hd__o21ai_4 c287 (.A1(net696),
    .A2(net708),
    .B1(net105),
    .Y(net789));
 sky130_fd_sc_hd__o21ai_2 c288 (.A1(net39),
    .A2(net12),
    .B1(net704),
    .Y(net122));
 sky130_fd_sc_hd__buf_4 c289 (.A(net606),
    .X(net790));
 sky130_fd_sc_hd__o21ai_4 c290 (.A1(net99),
    .A2(net861),
    .B1(net14),
    .Y(net820));
 sky130_fd_sc_hd__o21bai_4 c291 (.A1(net106),
    .A2(net869),
    .B1_N(net567),
    .Y(net123));
 sky130_fd_sc_hd__a21bo_4 c292 (.A1(net695),
    .A2(net29),
    .B1_N(net10),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 c293 (.A(net606),
    .X(net125));
 sky130_fd_sc_hd__sdfbbn_2 c294 (.CLK_N(clknet_4_2_0_clk),
    .D(net123),
    .RESET_B(net708),
    .SCD(net820),
    .SCE(net125),
    .SET_B(net891),
    .Q(net127),
    .Q_N(net126));
 sky130_fd_sc_hd__a21bo_1 c295 (.A1(net46),
    .A2(net124),
    .B1_N(net695),
    .X(net128));
 sky130_fd_sc_hd__a21o_1 c296 (.A1(net121),
    .A2(net46),
    .B1(net124),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 c297 (.A(net588),
    .X(net130));
 sky130_fd_sc_hd__a31oi_1 c298 (.A1(net124),
    .A2(net703),
    .A3(net130),
    .B1(net906),
    .Y(net131));
 sky130_fd_sc_hd__a41oi_1 c299 (.A1(net128),
    .A2(net124),
    .A3(net696),
    .A4(net131),
    .B1(net706),
    .Y(net132));
 sky130_fd_sc_hd__inv_1 c300 (.A(net588),
    .Y(net133));
 sky130_fd_sc_hd__a41o_1 c301 (.A1(net38),
    .A2(net130),
    .A3(net704),
    .A4(net790),
    .B1(net133),
    .X(net134));
 sky130_fd_sc_hd__sdfbbn_2 c302 (.CLK_N(clknet_4_2_0_clk),
    .D(net923),
    .RESET_B(net859),
    .SCD(net122),
    .SCE(net704),
    .SET_B(net128),
    .Q(net783),
    .Q_N(net135));
 sky130_fd_sc_hd__a41o_1 c303 (.A1(net134),
    .A2(net783),
    .A3(net789),
    .A4(net130),
    .B1(net607),
    .X(net136));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net136),
    .A1(net695),
    .A2(net133),
    .A3(net820),
    .S0(net134),
    .S1(net701),
    .X(net137));
 sky130_fd_sc_hd__o21ba_1 c305 (.A1(net131),
    .A2(net123),
    .B1_N(net130),
    .X(net138));
 sky130_fd_sc_hd__a21o_4 c306 (.A1(net138),
    .A2(net135),
    .B1(net606),
    .X(net787));
 sky130_fd_sc_hd__a41o_1 c307 (.A1(net708),
    .A2(net133),
    .A3(net135),
    .A4(net138),
    .B1(net607),
    .X(net139));
 sky130_fd_sc_hd__inv_1 c308 (.A(net605),
    .Y(net140));
 sky130_fd_sc_hd__a31o_4 c309 (.A1(net49),
    .A2(net870),
    .A3(net732),
    .B1(net31),
    .X(net141));
 sky130_fd_sc_hd__a21boi_4 c310 (.A1(net109),
    .A2(net736),
    .B1_N(net864),
    .Y(net142));
 sky130_fd_sc_hd__a31oi_4 c311 (.A1(net692),
    .A2(net109),
    .A3(net130),
    .B1(net141),
    .Y(net143));
 sky130_fd_sc_hd__xnor2_1 c312 (.A(net143),
    .B(net142),
    .Y(net144));
 sky130_fd_sc_hd__a31oi_1 c313 (.A1(net136),
    .A2(net30),
    .A3(net141),
    .B1(net567),
    .Y(net145));
 sky130_fd_sc_hd__a31o_4 c314 (.A1(net48),
    .A2(net735),
    .A3(net31),
    .B1(net692),
    .X(net146));
 sky130_fd_sc_hd__xor2_1 c315 (.A(net146),
    .B(net958),
    .X(net147));
 sky130_fd_sc_hd__o21bai_4 c316 (.A1(net130),
    .A2(net141),
    .B1_N(net146),
    .Y(net148));
 sky130_fd_sc_hd__xor2_4 c317 (.A(net142),
    .B(net143),
    .X(net149));
 sky130_fd_sc_hd__a21bo_1 c318 (.A1(net700),
    .A2(net903),
    .B1_N(net149),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 c319 (.A(net576),
    .X(net151));
 sky130_fd_sc_hd__mux2_4 c320 (.A0(net148),
    .A1(net140),
    .S(net151),
    .X(net815));
 sky130_fd_sc_hd__sdfbbp_1 c321 (.CLK(clknet_4_8_0_clk),
    .D(net150),
    .RESET_B(net151),
    .SCD(net147),
    .SCE(net149),
    .SET_B(net815),
    .Q(net784),
    .Q_N(net152));
 sky130_fd_sc_hd__clkbuf_2 c322 (.A(net605),
    .X(net153));
 sky130_fd_sc_hd__o21bai_2 c323 (.A1(net153),
    .A2(net144),
    .B1_N(net141),
    .Y(net154));
 sky130_fd_sc_hd__buf_6 c324 (.A(net539),
    .X(net155));
 sky130_fd_sc_hd__inv_6 c325 (.A(net539),
    .Y(net156));
 sky130_fd_sc_hd__a31oi_1 c326 (.A1(net151),
    .A2(net154),
    .A3(net882),
    .B1(net141),
    .Y(net157));
 sky130_fd_sc_hd__a31o_1 c327 (.A1(net952),
    .A2(net30),
    .A3(net882),
    .B1(net714),
    .X(net158));
 sky130_fd_sc_hd__a41o_1 c328 (.A1(net144),
    .A2(net151),
    .A3(net152),
    .A4(net130),
    .B1(net882),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net158),
    .A1(net154),
    .A2(net882),
    .A3(net153),
    .S0(net859),
    .S1(net146),
    .X(net160));
 sky130_fd_sc_hd__a31o_1 c330 (.A1(net76),
    .A2(net958),
    .A3(net155),
    .B1(net120),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 c331 (.A(net680),
    .X(net162));
 sky130_fd_sc_hd__a21bo_1 c332 (.A1(net790),
    .A2(net827),
    .B1_N(net606),
    .X(net163));
 sky130_fd_sc_hd__sdfbbn_1 c333 (.CLK_N(clknet_4_8_0_clk),
    .D(net762),
    .RESET_B(net73),
    .SCD(net887),
    .SCE(net884),
    .SET_B(net163),
    .Q(net165),
    .Q_N(net164));
 sky130_fd_sc_hd__a41oi_1 c334 (.A1(net159),
    .A2(net784),
    .A3(net73),
    .A4(net872),
    .B1(net921),
    .Y(net166));
 sky130_fd_sc_hd__o21bai_1 c335 (.A1(net73),
    .A2(net165),
    .B1_N(net800),
    .Y(net167));
 sky130_fd_sc_hd__inv_4 c336 (.A(net679),
    .Y(net168));
 sky130_fd_sc_hd__o21ba_2 c337 (.A1(net105),
    .A2(net870),
    .B1_N(net875),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(net168),
    .A1(net815),
    .A2(net832),
    .A3(net735),
    .S0(net875),
    .S1(net592),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 c339 (.A0(net169),
    .A1(net84),
    .A2(net762),
    .A3(net875),
    .S0(net591),
    .S1(net800),
    .X(net171));
 sky130_fd_sc_hd__a41oi_4 c340 (.A1(net169),
    .A2(net148),
    .A3(net876),
    .A4(net164),
    .B1(net560),
    .Y(net172));
 sky130_fd_sc_hd__a41o_1 c341 (.A1(net78),
    .A2(net875),
    .A3(net165),
    .A4(net887),
    .B1(net76),
    .X(net173));
 sky130_fd_sc_hd__a31o_4 c342 (.A1(net106),
    .A2(net865),
    .A3(net77),
    .B1(net875),
    .X(net848));
 sky130_fd_sc_hd__sdfbbn_1 c343 (.CLK_N(clknet_4_10_0_clk),
    .D(net169),
    .RESET_B(net159),
    .SCD(net172),
    .SCE(net875),
    .SET_B(net609),
    .Q(net175),
    .Q_N(net174));
 sky130_fd_sc_hd__mux4_2 c344 (.A0(net173),
    .A1(net168),
    .A2(net175),
    .A3(net148),
    .S0(net746),
    .S1(net848),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 c345 (.A(net574),
    .X(net177));
 sky130_fd_sc_hd__sdfbbp_1 c346 (.CLK(clknet_4_8_0_clk),
    .D(net162),
    .RESET_B(net176),
    .SCD(net77),
    .SCE(net820),
    .SET_B(net875),
    .Q(net179),
    .Q_N(net178));
 sky130_fd_sc_hd__a41oi_4 c347 (.A1(net148),
    .A2(net864),
    .A3(net178),
    .A4(net149),
    .B1(net876),
    .Y(net180));
 sky130_fd_sc_hd__mux4_2 c348 (.A0(net149),
    .A1(net179),
    .A2(net172),
    .A3(net177),
    .S0(net876),
    .S1(net604),
    .X(net824));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net176),
    .A1(net168),
    .A2(net180),
    .A3(net10),
    .S0(net178),
    .S1(net876),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net180),
    .A1(net914),
    .A2(net176),
    .A3(net875),
    .S0(net604),
    .S1(net613),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net177),
    .A1(net709),
    .A2(net176),
    .A3(net180),
    .S0(net560),
    .S1(net936),
    .X(net183));
 sky130_fd_sc_hd__a41o_1 c352 (.A1(net883),
    .A2(net882),
    .A3(net92),
    .A4(net877),
    .B1(net610),
    .X(net184));
 sky130_fd_sc_hd__a31o_1 c353 (.A1(net3),
    .A2(net746),
    .A3(net903),
    .B1(net877),
    .X(net830));
 sky130_fd_sc_hd__a31o_2 c354 (.A1(net870),
    .A2(net169),
    .A3(net94),
    .B1(net886),
    .X(net185));
 sky130_fd_sc_hd__a41o_1 c355 (.A1(net820),
    .A2(net93),
    .A3(net736),
    .A4(net609),
    .B1(net927),
    .X(net186));
 sky130_fd_sc_hd__mux4_2 c356 (.A0(net175),
    .A1(net778),
    .A2(net856),
    .A3(net755),
    .S0(net574),
    .S1(net611),
    .X(net808));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net165),
    .A1(net882),
    .A2(net808),
    .A3(net869),
    .S0(net180),
    .S1(net777),
    .X(net187));
 sky130_fd_sc_hd__mux4_4 c358 (.A0(net185),
    .A1(net718),
    .A2(net95),
    .A3(net777),
    .S0(net908),
    .S1(net824),
    .X(net188));
 sky130_fd_sc_hd__a31oi_4 c359 (.A1(net184),
    .A2(net827),
    .A3(net92),
    .B1(clknet_1_0__leaf_net616),
    .Y(net189));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net752),
    .A1(net789),
    .A2(net815),
    .A3(net164),
    .S0(net877),
    .S1(net777),
    .X(net190));
 sky130_fd_sc_hd__mux4_2 c361 (.A0(net881),
    .A1(net185),
    .A2(net808),
    .A3(net872),
    .S0(net828),
    .S1(net615),
    .X(net191));
 sky130_fd_sc_hd__mux4_2 c362 (.A0(net190),
    .A1(net778),
    .A2(net3),
    .A3(net823),
    .S0(net93),
    .S1(clknet_1_0__leaf_net616),
    .X(net192));
 sky130_fd_sc_hd__mux4_4 c363 (.A0(net191),
    .A1(net808),
    .A2(net877),
    .A3(net103),
    .S0(net828),
    .S1(clknet_1_0__leaf_net616),
    .X(net822));
 sky130_fd_sc_hd__a31oi_1 c364 (.A1(net866),
    .A2(net826),
    .A3(net184),
    .B1(clknet_1_0__leaf_net616),
    .Y(net834));
 sky130_fd_sc_hd__mux4_2 c365 (.A0(net92),
    .A1(net865),
    .A2(net91),
    .A3(net169),
    .S0(net3),
    .S1(net882),
    .X(net833));
 sky130_fd_sc_hd__mux4_1 c366 (.A0(net93),
    .A1(net827),
    .A2(net833),
    .A3(net830),
    .S0(net705),
    .S1(net609),
    .X(net193));
 sky130_fd_sc_hd__mux4_4 c367 (.A0(net180),
    .A1(net823),
    .A2(net874),
    .A3(net908),
    .S0(net777),
    .S1(net752),
    .X(net194));
 sky130_fd_sc_hd__mux4_4 c368 (.A0(net818),
    .A1(net848),
    .A2(net185),
    .A3(net609),
    .S0(clknet_1_1__leaf_net616),
    .S1(clknet_1_0__leaf_net617),
    .X(net195));
 sky130_fd_sc_hd__sdfbbn_1 c369 (.CLK_N(clknet_4_11_0_clk),
    .D(net190),
    .RESET_B(net93),
    .SCD(net705),
    .SCE(net778),
    .SET_B(clknet_1_0__leaf_net617),
    .Q(net197),
    .Q_N(net196));
 sky130_fd_sc_hd__mux4_4 c370 (.A0(net197),
    .A1(net883),
    .A2(net823),
    .A3(net886),
    .S0(net614),
    .S1(clknet_1_0__leaf_net803),
    .X(net198));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net88),
    .A1(net191),
    .A2(net833),
    .A3(net92),
    .S0(net818),
    .S1(net615),
    .X(net199));
 sky130_fd_sc_hd__mux4_2 c372 (.A0(clknet_1_0__leaf_net822),
    .A1(net196),
    .A2(net887),
    .A3(net828),
    .S0(net618),
    .S1(net620),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(clknet_1_0__leaf_net834),
    .A1(clknet_1_1__leaf_net200),
    .A2(net856),
    .A3(net3),
    .S0(clknet_1_1__leaf_net617),
    .S1(net619),
    .X(net807));
 sky130_fd_sc_hd__xor2_2 c396 (.A(net761),
    .B(net867),
    .X(net201));
 sky130_fd_sc_hd__xnor2_2 c397 (.A(net948),
    .B(net112),
    .Y(net202));
 sky130_fd_sc_hd__a21boi_2 c398 (.A1(net15),
    .A2(net690),
    .B1_N(net891),
    .Y(net203));
 sky130_fd_sc_hd__xnor2_4 c399 (.A(net11),
    .B(net880),
    .Y(net204));
 sky130_fd_sc_hd__mux2_1 c400 (.A0(net201),
    .A1(net761),
    .S(net891),
    .X(net205));
 sky130_fd_sc_hd__clkinv_8 c401 (.A(net561),
    .Y(net206));
 sky130_fd_sc_hd__o21bai_2 c402 (.A1(net685),
    .A2(net202),
    .B1_N(net206),
    .Y(net207));
 sky130_fd_sc_hd__o21bai_2 c403 (.A1(net202),
    .A2(net15),
    .B1_N(net206),
    .Y(net208));
 sky130_fd_sc_hd__o21a_4 c404 (.A1(net867),
    .A2(net207),
    .B1(net573),
    .X(net209));
 sky130_fd_sc_hd__xor2_2 c405 (.A(net203),
    .B(net201),
    .X(net210));
 sky130_fd_sc_hd__o21a_4 c406 (.A1(net209),
    .A2(net204),
    .B1(net761),
    .X(net211));
 sky130_fd_sc_hd__xnor2_2 c407 (.A(net209),
    .B(net573),
    .Y(net212));
 sky130_fd_sc_hd__a21o_1 c408 (.A1(net210),
    .A2(net868),
    .B1(net572),
    .X(net213));
 sky130_fd_sc_hd__mux4_2 c409 (.A0(net212),
    .A1(net108),
    .A2(net207),
    .A3(net209),
    .S0(net117),
    .S1(net211),
    .X(net214));
 sky130_fd_sc_hd__buf_4 c410 (.A(net561),
    .X(net215));
 sky130_fd_sc_hd__o21bai_2 c411 (.A1(net214),
    .A2(net215),
    .B1_N(net211),
    .Y(net216));
 sky130_fd_sc_hd__buf_4 c412 (.A(net561),
    .X(net217));
 sky130_fd_sc_hd__mux4_2 c413 (.A0(net203),
    .A1(net116),
    .A2(net205),
    .A3(net206),
    .S0(net214),
    .S1(net211),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net218),
    .A1(net203),
    .A2(net868),
    .A3(net215),
    .S0(net216),
    .S1(net211),
    .X(net219));
 sky130_fd_sc_hd__sdfbbn_1 c415 (.CLK_N(clknet_4_0_0_clk),
    .D(net217),
    .RESET_B(net103),
    .SCD(net216),
    .SCE(net110),
    .SET_B(net622),
    .Q(net221),
    .Q_N(net220));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net221),
    .A1(net217),
    .A2(net110),
    .A3(net215),
    .S0(net868),
    .S1(net218),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 c417 (.A(net561),
    .X(net223));
 sky130_fd_sc_hd__buf_6 c418 (.A(net589),
    .X(net224));
 sky130_fd_sc_hd__sdfbbp_1 c419 (.CLK(clknet_4_0_0_clk),
    .D(net207),
    .RESET_B(net210),
    .SCD(net714),
    .SCE(net129),
    .SET_B(net623),
    .Q(net226),
    .Q_N(net225));
 sky130_fd_sc_hd__buf_16 c420 (.A(net558),
    .X(net227));
 sky130_fd_sc_hd__a21o_1 c421 (.A1(net224),
    .A2(net909),
    .B1(net869),
    .X(net228));
 sky130_fd_sc_hd__o21bai_4 c422 (.A1(net206),
    .A2(net607),
    .B1_N(net623),
    .Y(net229));
 sky130_fd_sc_hd__o21bai_4 c423 (.A1(net704),
    .A2(net229),
    .B1_N(net123),
    .Y(net230));
 sky130_fd_sc_hd__xnor2_1 c424 (.A(net121),
    .B(net127),
    .Y(net231));
 sky130_fd_sc_hd__xor2_1 c425 (.A(net139),
    .B(net567),
    .X(net232));
 sky130_fd_sc_hd__inv_4 c426 (.A(net558),
    .Y(net233));
 sky130_fd_sc_hd__a31oi_2 c427 (.A1(net230),
    .A2(net210),
    .A3(net891),
    .B1(net622),
    .Y(net234));
 sky130_fd_sc_hd__a21boi_2 c428 (.A1(net231),
    .A2(net112),
    .B1_N(net121),
    .Y(net235));
 sky130_fd_sc_hd__xnor2_1 c429 (.A(net226),
    .B(net233),
    .Y(net236));
 sky130_fd_sc_hd__clkbuf_2 c430 (.A(net589),
    .X(net237));
 sky130_fd_sc_hd__o21ba_1 c431 (.A1(net236),
    .A2(net235),
    .B1_N(net228),
    .X(net238));
 sky130_fd_sc_hd__a31o_2 c432 (.A1(net40),
    .A2(net238),
    .A3(net235),
    .B1(net211),
    .X(net239));
 sky130_fd_sc_hd__mux2_2 c433 (.A0(net205),
    .A1(net139),
    .S(net225),
    .X(net240));
 sky130_fd_sc_hd__o21bai_4 c434 (.A1(net235),
    .A2(net228),
    .B1_N(net239),
    .Y(net821));
 sky130_fd_sc_hd__mux4_4 c435 (.A0(net237),
    .A1(net240),
    .A2(net714),
    .A3(net866),
    .S0(net208),
    .S1(net229),
    .X(net241));
 sky130_fd_sc_hd__a31o_1 c436 (.A1(net230),
    .A2(net229),
    .A3(net239),
    .B1(net624),
    .X(net242));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net238),
    .A1(net235),
    .A2(net236),
    .A3(net242),
    .S0(net139),
    .S1(net230),
    .X(net243));
 sky130_fd_sc_hd__a41oi_1 c438 (.A1(net228),
    .A2(net237),
    .A3(net238),
    .A4(net559),
    .B1(net624),
    .Y(net244));
 sky130_fd_sc_hd__clkbuf_2 c439 (.A(net593),
    .X(net245));
 sky130_fd_sc_hd__sdfrbp_1 c440 (.CLK(clknet_4_9_0_clk),
    .D(net240),
    .RESET_B(net141),
    .SCD(net8),
    .SCE(net204),
    .Q(net247),
    .Q_N(net246));
 sky130_fd_sc_hd__a21boi_2 c441 (.A1(net233),
    .A2(net239),
    .B1_N(net789),
    .Y(net248));
 sky130_fd_sc_hd__sdfrbp_1 c442 (.CLK(clknet_4_9_0_clk),
    .D(net248),
    .RESET_B(net861),
    .SCD(net869),
    .SCE(net882),
    .Q(net250),
    .Q_N(net249));
 sky130_fd_sc_hd__a21o_2 c443 (.A1(net247),
    .A2(net864),
    .B1(net239),
    .X(net251));
 sky130_fd_sc_hd__buf_1 c444 (.A(net588),
    .X(net252));
 sky130_fd_sc_hd__sdfrtn_1 c445 (.CLK_N(clknet_4_8_0_clk),
    .D(net30),
    .RESET_B(net910),
    .SCD(net251),
    .SCE(net858),
    .Q(net253));
 sky130_fd_sc_hd__sdfrtp_2 c446 (.CLK(clknet_4_2_0_clk),
    .D(net141),
    .RESET_B(net239),
    .SCD(net125),
    .SCE(net251),
    .Q(net254));
 sky130_fd_sc_hd__a41oi_4 c447 (.A1(net252),
    .A2(net253),
    .A3(net55),
    .A4(net254),
    .B1(net703),
    .Y(net255));
 sky130_fd_sc_hd__a41o_1 c448 (.A1(net254),
    .A2(net894),
    .A3(net237),
    .A4(net204),
    .B1(net623),
    .X(net256));
 sky130_fd_sc_hd__a31o_1 c449 (.A1(net204),
    .A2(net250),
    .A3(net725),
    .B1(net246),
    .X(net257));
 sky130_fd_sc_hd__buf_2 c450 (.A(net588),
    .X(net805));
 sky130_fd_sc_hd__sdfbbn_1 c451 (.CLK_N(clknet_4_9_0_clk),
    .D(net930),
    .RESET_B(net805),
    .SCD(net257),
    .SCE(net248),
    .SET_B(net935),
    .Q(net259),
    .Q_N(net258));
 sky130_fd_sc_hd__sdfrtp_2 c452 (.CLK(clknet_4_2_0_clk),
    .D(net252),
    .RESET_B(net248),
    .SCD(net259),
    .SCE(net894),
    .Q(net260));
 sky130_fd_sc_hd__sdfbbn_1 c453 (.CLK_N(clknet_4_9_0_clk),
    .D(net256),
    .RESET_B(net251),
    .SCD(net934),
    .SCE(net254),
    .SET_B(net260),
    .Q(net262),
    .Q_N(net261));
 sky130_fd_sc_hd__a41oi_1 c454 (.A1(net251),
    .A2(net209),
    .A3(net255),
    .A4(net253),
    .B1(net805),
    .Y(net263));
 sky130_fd_sc_hd__sdfbbp_1 c455 (.CLK(clknet_4_9_0_clk),
    .D(net140),
    .RESET_B(net253),
    .SCD(net256),
    .SCE(net240),
    .SET_B(net261),
    .Q(net793),
    .Q_N(net264));
 sky130_fd_sc_hd__sdfrtp_1 c456 (.CLK(clknet_4_3_0_clk),
    .D(net259),
    .RESET_B(net922),
    .SCD(net858),
    .SCE(net623),
    .Q(net265));
 sky130_fd_sc_hd__a31oi_2 c457 (.A1(net265),
    .A2(net706),
    .A3(net103),
    .B1(net264),
    .Y(net266));
 sky130_fd_sc_hd__a31oi_4 c458 (.A1(net793),
    .A2(net266),
    .A3(net255),
    .B1(net920),
    .Y(net802));
 sky130_fd_sc_hd__sdfbbn_1 c459 (.CLK_N(clknet_4_9_0_clk),
    .D(net257),
    .RESET_B(net150),
    .SCD(net265),
    .SCE(net125),
    .SET_B(net920),
    .Q(net268),
    .Q_N(net267));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net266),
    .A1(net260),
    .A2(net267),
    .A3(net787),
    .S0(net874),
    .S1(net255),
    .X(net269));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net256),
    .A1(net253),
    .A2(net269),
    .A3(net802),
    .S0(net268),
    .S1(net794),
    .X(net270));
 sky130_fd_sc_hd__o21ai_1 c462 (.A1(net884),
    .A2(net805),
    .B1(net760),
    .Y(net271));
 sky130_fd_sc_hd__o21ba_1 c463 (.A1(net760),
    .A2(net848),
    .B1_N(net718),
    .X(net272));
 sky130_fd_sc_hd__o21ba_1 c464 (.A1(net255),
    .A2(net272),
    .B1_N(net271),
    .X(net273));
 sky130_fd_sc_hd__o21ai_1 c465 (.A1(net768),
    .A2(net262),
    .B1(net227),
    .Y(net274));
 sky130_fd_sc_hd__a21bo_2 c466 (.A1(net272),
    .A2(net274),
    .B1_N(net172),
    .X(net785));
 sky130_fd_sc_hd__a31oi_2 c467 (.A1(net247),
    .A2(net703),
    .A3(net255),
    .B1(net887),
    .Y(net275));
 sky130_fd_sc_hd__o21a_1 c468 (.A1(net274),
    .A2(net227),
    .B1(net848),
    .X(net809));
 sky130_fd_sc_hd__a21bo_2 c469 (.A1(net273),
    .A2(net179),
    .B1_N(net275),
    .X(net799));
 sky130_fd_sc_hd__dlymetal6s2s_1 c470 (.A(net682),
    .X(net801));
 sky130_fd_sc_hd__inv_2 c471 (.A(net681),
    .Y(net276));
 sky130_fd_sc_hd__mux4_2 c472 (.A0(net275),
    .A1(net255),
    .A2(net77),
    .A3(net155),
    .S0(net168),
    .S1(net864),
    .X(net816));
 sky130_fd_sc_hd__a21o_1 c473 (.A1(net172),
    .A2(net815),
    .B1(net610),
    .X(net277));
 sky130_fd_sc_hd__sdfbbn_2 c474 (.CLK_N(clknet_4_11_0_clk),
    .D(net77),
    .RESET_B(net768),
    .SCD(net799),
    .SCE(net876),
    .SET_B(net918),
    .Q(net806),
    .Q_N(net278));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net179),
    .A1(net806),
    .A2(net275),
    .A3(net888),
    .S0(net816),
    .S1(net703),
    .X(net279));
 sky130_fd_sc_hd__a21boi_1 c476 (.A1(net31),
    .A2(net278),
    .B1_N(net77),
    .Y(net280));
 sky130_fd_sc_hd__buf_6 c477 (.A(net576),
    .X(net281));
 sky130_fd_sc_hd__a21bo_1 c478 (.A1(net276),
    .A2(net280),
    .B1_N(net279),
    .X(net282));
 sky130_fd_sc_hd__sdfbbp_1 c479 (.CLK(clknet_4_9_0_clk),
    .D(net262),
    .RESET_B(net279),
    .SCD(net282),
    .SCE(net77),
    .SET_B(net866),
    .Q(net284),
    .Q_N(net283));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net282),
    .A1(net284),
    .A2(net821),
    .A3(net882),
    .S0(net848),
    .S1(net77),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net168),
    .A1(net284),
    .A2(net172),
    .A3(net282),
    .S0(net865),
    .S1(net876),
    .X(net286));
 sky130_fd_sc_hd__a41o_1 c482 (.A1(net864),
    .A2(net271),
    .A3(net282),
    .A4(net276),
    .B1(net933),
    .X(net287));
 sky130_fd_sc_hd__sdfbbn_1 c483 (.CLK_N(clknet_4_9_0_clk),
    .D(net280),
    .RESET_B(net282),
    .SCD(net281),
    .SCE(net283),
    .SET_B(net563),
    .Q(net289),
    .Q_N(net288));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net725),
    .A1(net815),
    .A2(net185),
    .A3(net877),
    .S0(net810),
    .S1(net614),
    .X(net290));
 sky130_fd_sc_hd__sdfbbn_1 c485 (.CLK_N(clknet_4_11_0_clk),
    .D(clknet_1_0__leaf_net200),
    .RESET_B(net865),
    .SCD(net799),
    .SCE(net856),
    .SET_B(net614),
    .Q(net292),
    .Q_N(net291));
 sky130_fd_sc_hd__sdfbbp_1 c486 (.CLK(clknet_4_11_0_clk),
    .D(clknet_1_0__leaf_net189),
    .RESET_B(net95),
    .SCD(net778),
    .SCE(net894),
    .SET_B(net916),
    .Q(net294),
    .Q_N(net293));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net91),
    .A1(net778),
    .A2(net815),
    .A3(net209),
    .S0(net799),
    .S1(net610),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net705),
    .A1(net273),
    .A2(net815),
    .A3(net809),
    .S0(net725),
    .S1(net866),
    .X(net296));
 sky130_fd_sc_hd__a41o_1 c489 (.A1(net945),
    .A2(net818),
    .A3(net442),
    .A4(net877),
    .B1(net625),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net292),
    .A1(net926),
    .A2(net815),
    .A3(net873),
    .S0(net296),
    .S1(net882),
    .X(net298));
 sky130_fd_sc_hd__a41oi_4 c491 (.A1(net209),
    .A2(net725),
    .A3(clknet_1_1__leaf_net189),
    .A4(net291),
    .B1(net615),
    .Y(net299));
 sky130_fd_sc_hd__a31o_1 c492 (.A1(net815),
    .A2(net865),
    .A3(net614),
    .B1(net615),
    .X(net300));
 sky130_fd_sc_hd__mux4_2 c493 (.A0(net881),
    .A1(net209),
    .A2(net888),
    .A3(net800),
    .S0(net614),
    .S1(net625),
    .X(net811));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net103),
    .A1(net848),
    .A2(net894),
    .A3(net799),
    .S0(net615),
    .S1(clknet_1_0__leaf_net803),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net296),
    .A1(net804),
    .A2(net879),
    .A3(net811),
    .S0(net888),
    .S1(net626),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net156),
    .A1(net784),
    .A2(net811),
    .A3(clknet_1_0__leaf_net807),
    .S0(net290),
    .S1(net626),
    .X(net798));
 sky130_fd_sc_hd__mux4_4 c497 (.A0(net290),
    .A1(net292),
    .A2(clknet_1_1__leaf_net200),
    .A3(net886),
    .S0(net801),
    .S1(net787),
    .X(net303));
 sky130_fd_sc_hd__sdfbbn_1 c498 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net303),
    .RESET_B(net886),
    .SCD(net908),
    .SCE(net879),
    .SET_B(clknet_1_1__leaf_net803),
    .Q(net305),
    .Q_N(net304));
 sky130_fd_sc_hd__mux4_2 c499 (.A0(net778),
    .A1(net886),
    .A2(net304),
    .A3(net881),
    .S0(clknet_1_0__leaf_net200),
    .S1(net626),
    .X(net840));
 sky130_fd_sc_hd__sdfbbn_1 c500 (.CLK_N(clknet_4_14_0_clk),
    .D(net942),
    .RESET_B(net802),
    .SCD(clknet_1_0__leaf_net303),
    .SCE(net610),
    .SET_B(net924),
    .Q(net307),
    .Q_N(net306));
 sky130_fd_sc_hd__mux4_4 c501 (.A0(clknet_1_0__leaf_net798),
    .A1(net886),
    .A2(net91),
    .A3(net601),
    .S0(net626),
    .S1(net627),
    .X(net308));
 sky130_fd_sc_hd__mux4_2 c502 (.A0(net300),
    .A1(net305),
    .A2(net877),
    .A3(clknet_1_0__leaf_net840),
    .S0(net789),
    .S1(net626),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net291),
    .A1(net306),
    .A2(net305),
    .A3(net910),
    .S0(net865),
    .S1(net629),
    .X(net797));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net307),
    .A1(net281),
    .A2(net817),
    .A3(net209),
    .S0(net304),
    .S1(net626),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net95),
    .A1(net310),
    .A2(net797),
    .A3(net894),
    .S0(net304),
    .S1(net628),
    .X(net812));
 sky130_fd_sc_hd__o21ai_1 c528 (.A1(net223),
    .A2(net761),
    .B1(net206),
    .Y(net311));
 sky130_fd_sc_hd__a31o_4 c529 (.A1(net201),
    .A2(net10),
    .A3(net223),
    .B1(net108),
    .X(net312));
 sky130_fd_sc_hd__a21oi_4 c530 (.A1(net19),
    .A2(net206),
    .B1(net312),
    .Y(net313));
 sky130_fd_sc_hd__xnor2_4 c531 (.A(net690),
    .B(net868),
    .Y(net314));
 sky130_fd_sc_hd__xnor2_2 c532 (.A(net108),
    .B(net312),
    .Y(net315));
 sky130_fd_sc_hd__a31o_1 c533 (.A1(net210),
    .A2(net863),
    .A3(net761),
    .B1(net216),
    .X(net316));
 sky130_fd_sc_hd__xnor2_4 c534 (.A(net313),
    .B(net867),
    .Y(net317));
 sky130_fd_sc_hd__xnor2_1 c535 (.A(net312),
    .B(net317),
    .Y(net318));
 sky130_fd_sc_hd__a21o_1 c536 (.A1(net223),
    .A2(net718),
    .B1(net573),
    .X(net319));
 sky130_fd_sc_hd__sdfsbp_1 c537 (.CLK(clknet_4_1_0_clk),
    .D(net318),
    .SCD(net215),
    .SCE(net317),
    .SET_B(net863),
    .Q(net321),
    .Q_N(net320));
 sky130_fd_sc_hd__sdfsbp_2 c538 (.CLK(clknet_4_1_0_clk),
    .D(net116),
    .SCD(net319),
    .SCE(net206),
    .SET_B(net318),
    .Q(net323),
    .Q_N(net322));
 sky130_fd_sc_hd__a41o_1 c539 (.A1(net868),
    .A2(net108),
    .A3(net213),
    .A4(net322),
    .B1(net598),
    .X(net324));
 sky130_fd_sc_hd__a21boi_4 c540 (.A1(net311),
    .A2(net319),
    .B1_N(net324),
    .Y(net325));
 sky130_fd_sc_hd__a31o_1 c541 (.A1(net319),
    .A2(net313),
    .A3(net324),
    .B1(net321),
    .X(net326));
 sky130_fd_sc_hd__a41oi_4 c542 (.A1(net321),
    .A2(net866),
    .A3(net317),
    .A4(net863),
    .B1(net761),
    .Y(net327));
 sky130_fd_sc_hd__mux4_2 c543 (.A0(net314),
    .A1(net863),
    .A2(net326),
    .A3(net319),
    .S0(net312),
    .S1(net114),
    .X(net328));
 sky130_fd_sc_hd__sdfstp_2 c544 (.CLK(clknet_4_0_0_clk),
    .D(net326),
    .SCD(net319),
    .SCE(net937),
    .SET_B(net116),
    .Q(net329));
 sky130_fd_sc_hd__mux4_4 c545 (.A0(net867),
    .A1(net329),
    .A2(net220),
    .A3(net327),
    .S0(net314),
    .S1(net863),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(net324),
    .A1(net329),
    .A2(net220),
    .A3(net326),
    .S0(net572),
    .S1(net623),
    .X(net331));
 sky130_fd_sc_hd__a31oi_1 c547 (.A1(net690),
    .A2(net325),
    .A3(net312),
    .B1(net919),
    .Y(net332));
 sky130_fd_sc_hd__sdfstp_4 c548 (.CLK(clknet_4_1_0_clk),
    .D(net329),
    .SCD(net318),
    .SCE(net925),
    .SET_B(net586),
    .Q(net333));
 sky130_fd_sc_hd__a31o_1 c549 (.A1(net333),
    .A2(net329),
    .A3(net598),
    .B1(net632),
    .X(net334));
 sky130_fd_sc_hd__inv_12 c550 (.A(net581),
    .Y(net335));
 sky130_fd_sc_hd__a21oi_1 c551 (.A1(net229),
    .A2(net787),
    .B1(net237),
    .Y(net336));
 sky130_fd_sc_hd__o21ai_4 c552 (.A1(net124),
    .A2(net335),
    .B1(net114),
    .Y(net337));
 sky130_fd_sc_hd__xnor2_4 c553 (.A(net329),
    .B(net333),
    .Y(net338));
 sky130_fd_sc_hd__o21bai_4 c554 (.A1(net112),
    .A2(net871),
    .B1_N(net338),
    .Y(net339));
 sky130_fd_sc_hd__clkbuf_1 c555 (.A(net581),
    .X(net340));
 sky130_fd_sc_hd__inv_2 c556 (.A(net593),
    .Y(net341));
 sky130_fd_sc_hd__o21ba_1 c557 (.A1(net114),
    .A2(net224),
    .B1_N(net861),
    .X(net342));
 sky130_fd_sc_hd__a21boi_4 c558 (.A1(net245),
    .A2(net339),
    .B1_N(net716),
    .Y(net343));
 sky130_fd_sc_hd__o21ai_4 c559 (.A1(net335),
    .A2(net343),
    .B1(net559),
    .Y(net344));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net221),
    .A1(net343),
    .A2(net329),
    .A3(net115),
    .S0(net342),
    .S1(net340),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net226),
    .A1(net341),
    .A2(net343),
    .A3(net123),
    .S0(net718),
    .S1(net234),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_1 c562 (.A(net593),
    .X(net347));
 sky130_fd_sc_hd__xor2_4 c563 (.A(net343),
    .B(net29),
    .X(net348));
 sky130_fd_sc_hd__buf_2 c564 (.A(net593),
    .X(net349));
 sky130_fd_sc_hd__inv_2 c565 (.A(net928),
    .Y(net350));
 sky130_fd_sc_hd__sdfbbp_1 c566 (.CLK(clknet_4_1_0_clk),
    .D(net346),
    .RESET_B(net350),
    .SCD(net341),
    .SCE(net349),
    .SET_B(net929),
    .Q(net352),
    .Q_N(net351));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(net29),
    .A1(net349),
    .A2(net224),
    .A3(net863),
    .S0(net348),
    .S1(net351),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net340),
    .A1(net352),
    .A2(net341),
    .A3(net326),
    .S0(net859),
    .S1(net225),
    .X(net354));
 sky130_fd_sc_hd__buf_6 c569 (.A(clknet_1_0__leaf_net595),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(clknet_1_0__leaf_net355),
    .A1(net346),
    .A2(net353),
    .A3(net347),
    .S0(net348),
    .S1(net701),
    .X(net356));
 sky130_fd_sc_hd__mux4_2 c571 (.A0(net353),
    .A1(net348),
    .A2(net124),
    .A3(net341),
    .S0(net582),
    .S1(net634),
    .X(net357));
 sky130_fd_sc_hd__a41oi_4 c572 (.A1(net863),
    .A2(net790),
    .A3(net352),
    .A4(net115),
    .B1(net623),
    .Y(net358));
 sky130_fd_sc_hd__sdfbbn_1 c573 (.CLK_N(clknet_4_3_0_clk),
    .D(net206),
    .RESET_B(net930),
    .SCD(net327),
    .SCE(net566),
    .SET_B(net634),
    .Q(net360),
    .Q_N(net359));
 sky130_fd_sc_hd__a31o_4 c574 (.A1(net358),
    .A2(net322),
    .A3(net146),
    .B1(net623),
    .X(net361));
 sky130_fd_sc_hd__sdfbbn_1 c575 (.CLK_N(clknet_4_3_0_clk),
    .D(net347),
    .RESET_B(net314),
    .SCD(net863),
    .SCE(net135),
    .SET_B(net327),
    .Q(net363),
    .Q_N(net362));
 sky130_fd_sc_hd__a31oi_1 c576 (.A1(net861),
    .A2(net363),
    .A3(net211),
    .B1(net146),
    .Y(net364));
 sky130_fd_sc_hd__sdfbbp_1 c577 (.CLK(clknet_4_12_0_clk),
    .D(net269),
    .RESET_B(net253),
    .SCD(net41),
    .SCE(net623),
    .SET_B(net915),
    .Q(net366),
    .Q_N(net365));
 sky130_fd_sc_hd__a31oi_2 c578 (.A1(net115),
    .A2(net237),
    .A3(net19),
    .B1(net264),
    .Y(net367));
 sky130_fd_sc_hd__a31oi_4 c579 (.A1(net871),
    .A2(net146),
    .A3(net863),
    .B1(net623),
    .Y(net368));
 sky130_fd_sc_hd__a41o_1 c580 (.A1(net367),
    .A2(net339),
    .A3(net894),
    .A4(net368),
    .B1(net631),
    .X(net369));
 sky130_fd_sc_hd__a41oi_2 c581 (.A1(net364),
    .A2(net716),
    .A3(net366),
    .A4(net874),
    .B1(net315),
    .Y(net370));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net368),
    .A1(net363),
    .A2(net367),
    .A3(net314),
    .S0(net315),
    .S1(net369),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net336),
    .A1(net146),
    .A2(net251),
    .A3(net362),
    .S0(net314),
    .S1(net155),
    .X(net372));
 sky130_fd_sc_hd__mux4_4 c584 (.A0(net369),
    .A1(net251),
    .A2(net706),
    .A3(net361),
    .S0(net365),
    .S1(clknet_1_0__leaf_net635),
    .X(net373));
 sky130_fd_sc_hd__mux4_4 c585 (.A0(net19),
    .A1(net265),
    .A2(net891),
    .A3(net338),
    .S0(net369),
    .S1(clknet_1_0__leaf_net636),
    .X(net374));
 sky130_fd_sc_hd__a41oi_1 c586 (.A1(net360),
    .A2(net362),
    .A3(net152),
    .A4(net603),
    .B1(clknet_1_1__leaf_net636),
    .Y(net375));
 sky130_fd_sc_hd__mux4_4 c587 (.A0(net375),
    .A1(net362),
    .A2(net269),
    .A3(net368),
    .S0(clknet_1_0__leaf_net635),
    .S1(clknet_1_1__leaf_net636),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net366),
    .A1(net206),
    .A2(net267),
    .A3(net566),
    .S0(clknet_1_0__leaf_net636),
    .S1(clknet_1_0__leaf_net637),
    .X(net377));
 sky130_fd_sc_hd__mux4_4 c589 (.A0(clknet_1_0__leaf_net377),
    .A1(net881),
    .A2(net227),
    .A3(net368),
    .S0(clknet_1_1__leaf_net636),
    .S1(net638),
    .X(net378));
 sky130_fd_sc_hd__a41oi_1 c590 (.A1(net363),
    .A2(net358),
    .A3(net268),
    .A4(net718),
    .B1(net603),
    .Y(net379));
 sky130_fd_sc_hd__mux4_4 c591 (.A0(net706),
    .A1(clknet_1_0__leaf_net378),
    .A2(net367),
    .A3(net863),
    .S0(clknet_1_0__leaf_net637),
    .S1(net638),
    .X(net380));
 sky130_fd_sc_hd__mux4_4 c592 (.A0(net379),
    .A1(clknet_1_1__leaf_net377),
    .A2(clknet_1_0__leaf_net378),
    .A3(net582),
    .S0(net623),
    .S1(clknet_1_0__leaf_net636),
    .X(net381));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net368),
    .A1(net359),
    .A2(net379),
    .A3(net586),
    .S0(clknet_1_1__leaf_net636),
    .S1(net640),
    .X(net382));
 sky130_fd_sc_hd__a31oi_4 c594 (.A1(net344),
    .A2(net794),
    .A3(net896),
    .B1(clknet_1_1__leaf_net635),
    .Y(net383));
 sky130_fd_sc_hd__inv_1 c595 (.A(net589),
    .Y(net384));
 sky130_fd_sc_hd__a41oi_4 c596 (.A1(net155),
    .A2(net865),
    .A3(net227),
    .A4(net787),
    .B1(net283),
    .Y(net385));
 sky130_fd_sc_hd__a41oi_2 c597 (.A1(net10),
    .A2(net289),
    .A3(net894),
    .A4(net385),
    .B1(net267),
    .Y(net386));
 sky130_fd_sc_hd__a41oi_2 c598 (.A1(net357),
    .A2(net785),
    .A3(net709),
    .A4(net351),
    .B1(net176),
    .Y(net387));
 sky130_fd_sc_hd__sdfbbn_1 c599 (.CLK_N(clknet_4_12_0_clk),
    .D(net357),
    .RESET_B(net935),
    .SCD(net859),
    .SCE(net608),
    .SET_B(clknet_1_0__leaf_net635),
    .Q(net389),
    .Q_N(net388));
 sky130_fd_sc_hd__a41o_2 c600 (.A1(net155),
    .A2(net787),
    .A3(net152),
    .A4(net288),
    .B1(clknet_1_1__leaf_net635),
    .X(net390));
 sky130_fd_sc_hd__a41oi_4 c601 (.A1(net384),
    .A2(net804),
    .A3(net888),
    .A4(net155),
    .B1(net630),
    .Y(net391));
 sky130_fd_sc_hd__mux4_2 c602 (.A0(net227),
    .A1(clknet_1_0__leaf_net355),
    .A2(net284),
    .A3(net804),
    .S0(net881),
    .S1(net264),
    .X(net392));
 sky130_fd_sc_hd__a41oi_4 c603 (.A1(net391),
    .A2(net317),
    .A3(net894),
    .A4(net804),
    .B1(clknet_1_1__leaf_net637),
    .Y(net393));
 sky130_fd_sc_hd__sdfbbn_1 c604 (.CLK_N(clknet_4_9_0_clk),
    .D(net277),
    .RESET_B(net289),
    .SCD(net865),
    .SCE(clknet_1_0__leaf_net393),
    .SET_B(clknet_1_1__leaf_net637),
    .Q(net395),
    .Q_N(net394));
 sky130_fd_sc_hd__sdfbbp_1 c605 (.CLK(clknet_4_12_0_clk),
    .D(net931),
    .RESET_B(net385),
    .SCD(net327),
    .SCE(net394),
    .SET_B(net859),
    .Q(net397),
    .Q_N(net396));
 sky130_fd_sc_hd__mux4_4 c606 (.A0(net268),
    .A1(net249),
    .A2(net881),
    .A3(clknet_1_1__leaf_net393),
    .S0(clknet_1_1__leaf_net355),
    .S1(net865),
    .X(net398));
 sky130_fd_sc_hd__a41o_2 c607 (.A1(net392),
    .A2(net389),
    .A3(net317),
    .A4(net396),
    .B1(net631),
    .X(net399));
 sky130_fd_sc_hd__a41oi_4 c608 (.A1(net390),
    .A2(net176),
    .A3(net397),
    .A4(clknet_1_0__leaf_net393),
    .B1(net848),
    .Y(net400));
 sky130_fd_sc_hd__mux4_2 c609 (.A0(net317),
    .A1(net396),
    .A2(clknet_1_0__leaf_net393),
    .A3(net395),
    .S0(clknet_1_0__leaf_net399),
    .S1(net608),
    .X(net401));
 sky130_fd_sc_hd__mux4_4 c610 (.A0(clknet_1_1__leaf_net399),
    .A1(net155),
    .A2(net176),
    .A3(net385),
    .S0(net388),
    .S1(net644),
    .X(net402));
 sky130_fd_sc_hd__a41o_2 c611 (.A1(net383),
    .A2(clknet_1_1__leaf_net393),
    .A3(net397),
    .A4(clknet_1_0__leaf_net378),
    .B1(net645),
    .X(net403));
 sky130_fd_sc_hd__mux4_4 c612 (.A0(net888),
    .A1(net866),
    .A2(clknet_1_1__leaf_net635),
    .A3(clknet_1_1__leaf_net637),
    .S0(net641),
    .S1(net644),
    .X(net404));
 sky130_fd_sc_hd__mux4_4 c613 (.A0(net395),
    .A1(clknet_1_1__leaf_net393),
    .A2(net264),
    .A3(net866),
    .S0(net814),
    .S1(net644),
    .X(net405));
 sky130_fd_sc_hd__mux4_2 c614 (.A0(net10),
    .A1(net804),
    .A2(clknet_1_0__leaf_net404),
    .A3(net590),
    .S0(net644),
    .S1(net645),
    .X(net406));
 sky130_fd_sc_hd__mux4_2 c615 (.A0(net406),
    .A1(clknet_1_0__leaf_net404),
    .A2(net603),
    .A3(net791),
    .S0(net644),
    .S1(net645),
    .X(net792));
 sky130_fd_sc_hd__mux4_4 c616 (.A0(net894),
    .A1(net804),
    .A2(net361),
    .A3(net211),
    .S0(net152),
    .S1(clknet_1_1__leaf_net840),
    .X(net407));
 sky130_fd_sc_hd__mux4_4 c617 (.A0(clknet_1_1__leaf_net309),
    .A1(clknet_1_0__leaf_net840),
    .A2(net185),
    .A3(net789),
    .S0(net327),
    .S1(net94),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net94),
    .A1(net185),
    .A2(net894),
    .A3(net304),
    .S0(net627),
    .S1(net649),
    .X(net409));
 sky130_fd_sc_hd__mux4_2 c619 (.A0(net785),
    .A1(clknet_1_1__leaf_net378),
    .A2(net784),
    .A3(net703),
    .S0(net879),
    .S1(net647),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net409),
    .A1(net873),
    .A2(net787),
    .A3(net793),
    .S0(net337),
    .S1(net630),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net337),
    .A1(net305),
    .A2(net91),
    .A3(net627),
    .S0(net640),
    .S1(net644),
    .X(net412));
 sky130_fd_sc_hd__mux4_4 c622 (.A0(net385),
    .A1(net886),
    .A2(net273),
    .A3(clknet_1_0__leaf_net309),
    .S0(net789),
    .S1(net650),
    .X(net413));
 sky130_fd_sc_hd__mux4_2 c623 (.A0(net273),
    .A1(net784),
    .A2(net211),
    .A3(net770),
    .S0(net865),
    .S1(net649),
    .X(net796));
 sky130_fd_sc_hd__mux4_2 c624 (.A0(net305),
    .A1(net804),
    .A2(net814),
    .A3(net135),
    .S0(net631),
    .S1(net652),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net211),
    .A1(net414),
    .A2(clknet_1_1__leaf_net378),
    .A3(net888),
    .S0(net627),
    .S1(net653),
    .X(net415));
 sky130_fd_sc_hd__mux4_2 c626 (.A0(net338),
    .A1(net881),
    .A2(net785),
    .A3(net793),
    .S0(net648),
    .S1(net653),
    .X(net829));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net327),
    .A1(net337),
    .A2(net94),
    .A3(net620),
    .S0(net641),
    .S1(net654),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net211),
    .A1(net888),
    .A2(net804),
    .A3(net648),
    .S0(net653),
    .S1(net654),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net397),
    .A1(net417),
    .A2(net91),
    .A3(net893),
    .S0(net649),
    .S1(clknet_1_0__leaf_net655),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net185),
    .A1(net794),
    .A2(net562),
    .A3(net646),
    .S0(net653),
    .S1(clknet_1_1__leaf_net655),
    .X(net419));
 sky130_fd_sc_hd__mux4_2 c631 (.A0(net414),
    .A1(net796),
    .A2(net648),
    .A3(net652),
    .S0(net653),
    .S1(clknet_1_1__leaf_net655),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(clknet_1_1__leaf_net378),
    .A1(net120),
    .A2(net796),
    .A3(net651),
    .S0(net653),
    .S1(net654),
    .X(net421));
 sky130_fd_sc_hd__mux4_2 c633 (.A0(net419),
    .A1(net414),
    .A2(net562),
    .A3(net619),
    .S0(net647),
    .S1(clknet_1_1__leaf_net656),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net770),
    .A1(net264),
    .A2(net651),
    .A3(net652),
    .S0(net654),
    .S1(clknet_1_1__leaf_net656),
    .X(net836));
 sky130_fd_sc_hd__mux4_4 c635 (.A0(clknet_1_1__leaf_net418),
    .A1(net152),
    .A2(net608),
    .A3(net652),
    .S0(clknet_1_0__leaf_net655),
    .S1(clknet_1_0__leaf_net656),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(clknet_1_1__leaf_net423),
    .A1(net829),
    .A2(net649),
    .A3(net650),
    .S0(clknet_1_0__leaf_net655),
    .S1(clknet_1_0__leaf_net656),
    .X(net424));
 sky130_fd_sc_hd__mux4_2 c637 (.A0(clknet_1_0__leaf_net423),
    .A1(net821),
    .A2(net414),
    .A3(clknet_1_0__leaf_net418),
    .S0(net590),
    .S1(net603),
    .X(net425));
 sky130_fd_sc_hd__xnor2_1 c660 (.A(net334),
    .B(net212),
    .Y(net426));
 sky130_fd_sc_hd__xor2_2 c661 (.A(net113),
    .B(net862),
    .X(net427));
 sky130_fd_sc_hd__xnor2_4 c662 (.A(net217),
    .B(net862),
    .Y(net428));
 sky130_fd_sc_hd__xor2_4 c663 (.A(net117),
    .B(net788),
    .X(net429));
 sky130_fd_sc_hd__o21a_1 c664 (.A1(net761),
    .A2(net428),
    .B1(net322),
    .X(net430));
 sky130_fd_sc_hd__xor2_1 c665 (.A(net110),
    .B(net427),
    .X(net431));
 sky130_fd_sc_hd__mux2_1 c666 (.A0(net113),
    .A1(net862),
    .S(net428),
    .X(net432));
 sky130_fd_sc_hd__sdfstp_1 c667 (.CLK(clknet_4_5_0_clk),
    .D(net427),
    .SCD(net325),
    .SCE(net862),
    .SET_B(net959),
    .Q(net433));
 sky130_fd_sc_hd__xnor2_1 c668 (.A(net212),
    .B(net433),
    .Y(net434));
 sky130_fd_sc_hd__buf_1 c669 (.A(net585),
    .X(net435));
 sky130_fd_sc_hd__a41o_1 c670 (.A1(net857),
    .A2(net334),
    .A3(net428),
    .A4(net862),
    .B1(net919),
    .X(net436));
 sky130_fd_sc_hd__mux2_1 c671 (.A0(net427),
    .A1(net862),
    .S(net585),
    .X(net437));
 sky130_fd_sc_hd__o21bai_2 c672 (.A1(net435),
    .A2(net862),
    .B1_N(net585),
    .Y(net438));
 sky130_fd_sc_hd__xor2_2 c673 (.A(net860),
    .B(net943),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c674 (.A0(net438),
    .A1(net428),
    .A2(net761),
    .A3(net437),
    .S0(net857),
    .S1(net862),
    .X(net440));
 sky130_fd_sc_hd__inv_4 c675 (.A(net585),
    .Y(net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__xnor2_1 c677 (.A(net428),
    .B(net860),
    .Y(net443));
 sky130_fd_sc_hd__mux2_1 c678 (.A0(net215),
    .A1(net438),
    .S(net427),
    .X(net444));
 sky130_fd_sc_hd__buf_1 c679 (.A(net684),
    .X(net445));
 sky130_fd_sc_hd__mux4_4 c680 (.A0(net441),
    .A1(net428),
    .A2(net443),
    .A3(net857),
    .S0(net438),
    .S1(net445),
    .X(net446));
 sky130_fd_sc_hd__o21ai_2 c681 (.A1(net445),
    .A2(net435),
    .B1(net660),
    .Y(net447));
 sky130_fd_sc_hd__a21bo_1 c682 (.A1(net335),
    .A2(net794),
    .B1_N(net123),
    .X(net448));
 sky130_fd_sc_hd__a31oi_1 c683 (.A1(net433),
    .A2(net333),
    .A3(net325),
    .B1(net660),
    .Y(net449));
 sky130_fd_sc_hd__sedfxbp_2 c684 (.CLK(clknet_4_4_0_clk),
    .D(net123),
    .DE(net448),
    .SCD(net862),
    .SCE(net659),
    .Q(net451),
    .Q_N(net450));
 sky130_fd_sc_hd__sedfxbp_1 c685 (.CLK(clknet_4_5_0_clk),
    .D(net862),
    .DE(net325),
    .SCD(net434),
    .SCE(net351),
    .Q(net453),
    .Q_N(net452));
 sky130_fd_sc_hd__clkbuf_2 c686 (.A(net541),
    .X(net454));
 sky130_fd_sc_hd__mux2_1 c687 (.A0(net453),
    .A1(net790),
    .S(net450),
    .X(net455));
 sky130_fd_sc_hd__sdfbbn_2 c688 (.CLK_N(clknet_4_4_0_clk),
    .D(net434),
    .RESET_B(net451),
    .SCD(net426),
    .SCE(net431),
    .SET_B(net455),
    .Q(net457),
    .Q_N(net456));
 sky130_fd_sc_hd__clkbuf_2 c689 (.A(net540),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net213),
    .A1(net230),
    .A2(net339),
    .A3(net348),
    .S0(net458),
    .S1(net660),
    .X(net459));
 sky130_fd_sc_hd__a41o_1 c691 (.A1(net457),
    .A2(net458),
    .A3(net230),
    .A4(net454),
    .B1(net860),
    .X(net460));
 sky130_fd_sc_hd__sdfbbn_1 c692 (.CLK_N(clknet_4_5_0_clk),
    .D(net458),
    .RESET_B(net460),
    .SCD(net339),
    .SCE(net135),
    .SET_B(net857),
    .Q(net462),
    .Q_N(net461));
 sky130_fd_sc_hd__a41o_1 c693 (.A1(net325),
    .A2(net458),
    .A3(net454),
    .A4(net860),
    .B1(net941),
    .X(net463));
 sky130_fd_sc_hd__sedfxtp_2 c694 (.CLK(clknet_4_5_0_clk),
    .D(net459),
    .DE(net448),
    .SCD(net455),
    .SCE(net860),
    .Q(net464));
 sky130_fd_sc_hd__a31o_1 c695 (.A1(net123),
    .A2(net464),
    .A3(net456),
    .B1(net624),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net234),
    .A1(net464),
    .A2(net857),
    .A3(net457),
    .S0(net448),
    .S1(net465),
    .X(net466));
 sky130_fd_sc_hd__a41o_2 c697 (.A1(net465),
    .A2(net458),
    .A3(net452),
    .A4(net583),
    .B1(net662),
    .X(net467));
 sky130_fd_sc_hd__mux4_4 c698 (.A0(net343),
    .A1(net352),
    .A2(net464),
    .A3(net333),
    .S0(net444),
    .S1(net584),
    .X(net468));
 sky130_fd_sc_hd__a41o_1 c699 (.A1(net224),
    .A2(net857),
    .A3(net349),
    .A4(net860),
    .B1(net913),
    .X(net469));
 sky130_fd_sc_hd__mux4_4 c700 (.A0(net430),
    .A1(net464),
    .A2(net461),
    .A3(net860),
    .S0(net624),
    .S1(net634),
    .X(net470));
 sky130_fd_sc_hd__a41o_1 c701 (.A1(net431),
    .A2(net230),
    .A3(net857),
    .A4(net597),
    .B1(net665),
    .X(net471));
 sky130_fd_sc_hd__mux4_2 c702 (.A0(net339),
    .A1(net453),
    .A2(net467),
    .A3(clknet_1_0__leaf_net595),
    .S0(net664),
    .S1(net665),
    .X(net472));
 sky130_fd_sc_hd__sedfxtp_2 c703 (.CLK(clknet_4_6_0_clk),
    .D(net348),
    .DE(clknet_1_0__leaf_net472),
    .SCD(net461),
    .SCE(net467),
    .Q(net473));
 sky130_fd_sc_hd__sedfxtp_4 c704 (.CLK(clknet_4_7_0_clk),
    .D(net447),
    .DE(net361),
    .SCD(net938),
    .SCE(net939),
    .Q(net474));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net454),
    .A1(net857),
    .A2(net462),
    .A3(net455),
    .S0(net467),
    .S1(net566),
    .X(net475));
 sky130_fd_sc_hd__a31o_1 c706 (.A1(net339),
    .A2(net451),
    .A3(net660),
    .B1(net666),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net447),
    .A1(net349),
    .A2(net339),
    .A3(net467),
    .S0(net454),
    .S1(net794),
    .X(net477));
 sky130_fd_sc_hd__sdfrbp_2 c708 (.CLK(clknet_4_6_0_clk),
    .D(net125),
    .RESET_B(clknet_1_1__leaf_net472),
    .SCD(net860),
    .SCE(net339),
    .Q(net479),
    .Q_N(net478));
 sky130_fd_sc_hd__mux4_2 c709 (.A0(net476),
    .A1(net899),
    .A2(net474),
    .A3(net868),
    .S0(net349),
    .S1(net478),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net439),
    .A1(net260),
    .A2(net447),
    .A3(net478),
    .S0(net873),
    .S1(net639),
    .X(net481));
 sky130_fd_sc_hd__mux4_4 c711 (.A0(net439),
    .A1(net467),
    .A2(net474),
    .A3(net478),
    .S0(net642),
    .S1(net885),
    .X(net482));
 sky130_fd_sc_hd__mux4_2 c712 (.A0(net260),
    .A1(net480),
    .A2(net454),
    .A3(net429),
    .S0(net633),
    .S1(net885),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net868),
    .A1(net323),
    .A2(net859),
    .A3(net640),
    .S0(net885),
    .S1(net932),
    .X(net484));
 sky130_fd_sc_hd__mux4_4 c714 (.A0(net898),
    .A1(net467),
    .A2(net361),
    .A3(net478),
    .S0(net633),
    .S1(net885),
    .X(net485));
 sky130_fd_sc_hd__mux4_2 c715 (.A0(net860),
    .A1(net127),
    .A2(net633),
    .A3(net639),
    .S0(net885),
    .S1(net932),
    .X(net486));
 sky130_fd_sc_hd__mux4_2 c716 (.A0(net873),
    .A1(net479),
    .A2(net456),
    .A3(net557),
    .S0(net624),
    .S1(net885),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(clknet_1_0__leaf_net483),
    .A1(net897),
    .A2(net486),
    .A3(net478),
    .S0(net938),
    .S1(net915),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net455),
    .A1(net783),
    .A2(net633),
    .A3(net666),
    .S0(net885),
    .S1(net669),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net55),
    .A1(net486),
    .A2(net868),
    .A3(clknet_1_1__leaf_net483),
    .S0(net566),
    .S1(net885),
    .X(net490));
 sky130_fd_sc_hd__mux4_4 c720 (.A0(net486),
    .A1(net429),
    .A2(net323),
    .A3(net473),
    .S0(net474),
    .S1(net671),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net474),
    .A1(net860),
    .A2(net857),
    .A3(net639),
    .S0(net940),
    .S1(net673),
    .X(net492));
 sky130_fd_sc_hd__mux4_2 c722 (.A0(net462),
    .A1(net873),
    .A2(net868),
    .A3(net624),
    .S0(net642),
    .S1(net673),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net489),
    .A1(net477),
    .A2(net479),
    .A3(net873),
    .S0(net493),
    .S1(net944),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net432),
    .A1(net479),
    .A2(net486),
    .A3(net556),
    .S0(net673),
    .S1(net946),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net457),
    .A1(net454),
    .A2(net493),
    .A3(clknet_1_0__leaf_net594),
    .S0(net643),
    .S1(net885),
    .X(net496));
 sky130_fd_sc_hd__mux4_2 c726 (.A0(net224),
    .A1(clknet_1_1__leaf_net496),
    .A2(net284),
    .A3(net487),
    .S0(net718),
    .S1(net661),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net703),
    .A1(net709),
    .A2(net461),
    .A3(net473),
    .S0(net878),
    .S1(net641),
    .X(net498));
 sky130_fd_sc_hd__mux4_4 c728 (.A0(net352),
    .A1(net473),
    .A2(clknet_1_0__leaf_net496),
    .A3(net479),
    .S0(net878),
    .S1(net640),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net323),
    .A1(net473),
    .A2(net478),
    .A3(net790),
    .S0(net661),
    .S1(net664),
    .X(net500));
 sky130_fd_sc_hd__mux4_2 c730 (.A0(net881),
    .A1(net451),
    .A2(net878),
    .A3(clknet_1_0__leaf_net499),
    .S0(net661),
    .S1(net664),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net462),
    .A1(net716),
    .A2(net866),
    .A3(net493),
    .S0(net487),
    .S1(net645),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net859),
    .A1(net896),
    .A2(net597),
    .A3(net645),
    .S0(net646),
    .S1(net664),
    .X(net503));
 sky130_fd_sc_hd__mux4_2 c733 (.A0(net479),
    .A1(clknet_1_0__leaf_net497),
    .A2(net896),
    .A3(net893),
    .S0(net661),
    .S1(net675),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net498),
    .A1(net479),
    .A2(clknet_1_0__leaf_net496),
    .A3(net716),
    .S0(net670),
    .S1(net675),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net487),
    .A1(net352),
    .A2(net878),
    .A3(net660),
    .S0(net885),
    .S1(net675),
    .X(net506));
 sky130_fd_sc_hd__mux4_2 c736 (.A0(net506),
    .A1(net284),
    .A2(clknet_1_0__leaf_net504),
    .A3(clknet_1_0__leaf_net505),
    .S0(clknet_1_0__leaf_net497),
    .S1(net660),
    .X(net507));
 sky130_fd_sc_hd__mux4_4 c737 (.A0(net127),
    .A1(clknet_1_0__leaf_net505),
    .A2(net456),
    .A3(clknet_1_0__leaf_net497),
    .S0(clknet_1_0__leaf_net504),
    .S1(net661),
    .X(net508));
 sky130_fd_sc_hd__mux4_4 c738 (.A0(net500),
    .A1(net501),
    .A2(net479),
    .A3(net224),
    .S0(net859),
    .S1(net645),
    .X(net509));
 sky130_fd_sc_hd__mux4_2 c739 (.A0(net893),
    .A1(net457),
    .A2(net878),
    .A3(net661),
    .S0(net669),
    .S1(clknet_1_0__leaf_net676),
    .X(net510));
 sky130_fd_sc_hd__mux4_2 c740 (.A0(net502),
    .A1(net493),
    .A2(net284),
    .A3(net878),
    .S0(clknet_1_0__leaf_net497),
    .S1(net661),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net510),
    .A1(net511),
    .A2(net127),
    .A3(net878),
    .S0(clknet_1_1__leaf_net505),
    .S1(net893),
    .X(net512));
 sky130_fd_sc_hd__mux4_2 c742 (.A0(clknet_1_1__leaf_net504),
    .A1(net783),
    .A2(net790),
    .A3(clknet_1_1__leaf_net404),
    .S0(net645),
    .S1(net660),
    .X(net513));
 sky130_fd_sc_hd__mux4_4 c743 (.A0(net512),
    .A1(net507),
    .A2(net866),
    .A3(clknet_1_0__leaf_net513),
    .S0(net896),
    .S1(net660),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net514),
    .A1(clknet_1_0__leaf_net513),
    .A2(net323),
    .A3(clknet_1_1__leaf_net504),
    .S0(net709),
    .S1(net661),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(clknet_1_1__leaf_net513),
    .A1(clknet_1_1__leaf_net497),
    .A2(net896),
    .A3(net351),
    .S0(net224),
    .S1(net578),
    .X(net516));
 sky130_fd_sc_hd__mux4_2 c746 (.A0(net508),
    .A1(net284),
    .A2(net873),
    .A3(net645),
    .S0(net661),
    .S1(net675),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net516),
    .A1(clknet_1_0__leaf_net517),
    .A2(net462),
    .A3(clknet_1_1__leaf_net513),
    .S0(net645),
    .S1(net670),
    .X(net518));
 sky130_fd_sc_hd__mux4_2 c748 (.A0(net94),
    .A1(clknet_1_0__leaf_net404),
    .A2(net701),
    .A3(net873),
    .S0(net646),
    .S1(clknet_1_1__leaf_net676),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net361),
    .A1(clknet_1_1__leaf_net404),
    .A2(net783),
    .A3(net577),
    .S0(net654),
    .S1(clknet_1_0__leaf_net676),
    .X(net520));
 sky130_fd_sc_hd__mux4_2 c750 (.A0(clknet_1_1__leaf_net404),
    .A1(net493),
    .A2(net879),
    .A3(clknet_1_0__leaf_net657),
    .S0(net667),
    .S1(clknet_1_0__leaf_net677),
    .X(net521));
 sky130_fd_sc_hd__mux4_4 c751 (.A0(net91),
    .A1(clknet_1_0__leaf_net521),
    .A2(net361),
    .A3(clknet_1_0__leaf_net404),
    .S0(net646),
    .S1(clknet_1_0__leaf_net677),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net361),
    .A1(clknet_1_0__leaf_net521),
    .A2(net91),
    .A3(net578),
    .S0(clknet_1_1__leaf_net657),
    .S1(net667),
    .X(net523));
 sky130_fd_sc_hd__mux4_4 c753 (.A0(net718),
    .A1(clknet_1_1__leaf_net521),
    .A2(clknet_1_1__leaf_net517),
    .A3(net567),
    .S0(clknet_1_1__leaf_net596),
    .S1(net654),
    .X(net524));
 sky130_fd_sc_hd__mux4_2 c754 (.A0(net519),
    .A1(clknet_1_0__leaf_net521),
    .A2(clknet_1_1__leaf_net404),
    .A3(net493),
    .S0(net654),
    .S1(net667),
    .X(net525));
 sky130_fd_sc_hd__mux4_2 c755 (.A0(net493),
    .A1(clknet_1_1__leaf_net497),
    .A2(clknet_1_0__leaf_net521),
    .A3(net878),
    .S0(net646),
    .S1(clknet_1_1__leaf_net677),
    .X(net526));
 sky130_fd_sc_hd__mux4_4 c756 (.A0(net525),
    .A1(clknet_1_0__leaf_net517),
    .A2(clknet_1_0__leaf_net526),
    .A3(net94),
    .S0(clknet_1_0__leaf_net521),
    .S1(clknet_1_1__leaf_net677),
    .X(net527));
 sky130_fd_sc_hd__mux4_4 c757 (.A0(net120),
    .A1(net493),
    .A2(clknet_1_0__leaf_net521),
    .A3(net646),
    .S0(clknet_1_0__leaf_net657),
    .S1(clknet_1_0__leaf_net677),
    .X(net528));
 sky130_fd_sc_hd__mux4_2 c758 (.A0(net878),
    .A1(clknet_1_1__leaf_net526),
    .A2(clknet_1_1__leaf_net521),
    .A3(clknet_1_1__leaf_net497),
    .S0(net577),
    .S1(clknet_1_1__leaf_net657),
    .X(net529));
 sky130_fd_sc_hd__mux4_2 c759 (.A0(clknet_1_1__leaf_net521),
    .A1(clknet_1_1__leaf_net517),
    .A2(net493),
    .A3(clknet_1_0__leaf_net596),
    .S0(net602),
    .S1(clknet_1_1__leaf_net677),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net716),
    .A1(clknet_1_1__leaf_net521),
    .A2(net878),
    .A3(net600),
    .S0(clknet_1_1__leaf_net676),
    .S1(clknet_1_0__leaf_net678),
    .X(net531));
 sky130_fd_sc_hd__mux4_2 c761 (.A0(net529),
    .A1(net531),
    .A2(clknet_1_1__leaf_net517),
    .A3(clknet_1_1__leaf_net404),
    .S0(net602),
    .S1(clknet_1_1__leaf_net678),
    .X(net532));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(clknet_1_1__leaf_net499),
    .A1(net795),
    .A2(clknet_1_1__leaf_net594),
    .A3(net641),
    .S0(clknet_1_0__leaf_net657),
    .S1(clknet_1_0__leaf_net678),
    .X(net533));
 sky130_fd_sc_hd__a41oi_1 merge763 (.A1(net216),
    .A2(net794),
    .A3(net238),
    .A4(net706),
    .B1(net821),
    .Y(net534));
 sky130_fd_sc_hd__mux4_1 merge764 (.A0(net858),
    .A1(net84),
    .A2(net875),
    .A3(net904),
    .S0(net576),
    .S1(net591),
    .X(net535));
 sky130_fd_sc_hd__a41oi_1 merge765 (.A1(net430),
    .A2(net434),
    .A3(net334),
    .A4(net857),
    .B1(net439),
    .Y(net536));
 sky130_fd_sc_hd__a41o_1 merge766 (.A1(net205),
    .A2(net120),
    .A3(net19),
    .A4(net202),
    .B1(net209),
    .X(net537));
 sky130_fd_sc_hd__a41oi_2 merge767 (.A1(net47),
    .A2(net106),
    .A3(net114),
    .A4(net36),
    .B1(net124),
    .Y(net538));
 sky130_fd_sc_hd__inv_4 merge768 (.A(net589),
    .Y(net539));
 sky130_fd_sc_hd__sdfrbp_1 merge769 (.CLK(clknet_4_5_0_clk),
    .D(net450),
    .RESET_B(net911),
    .SCD(net444),
    .SCE(net456),
    .Q(net541),
    .Q_N(net540));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(net858),
    .A1(net77),
    .A2(net103),
    .A3(net799),
    .S0(net895),
    .S1(net579),
    .X(net542));
 sky130_fd_sc_hd__a41oi_1 merge771 (.A1(net236),
    .A2(net209),
    .A3(net251),
    .A4(net239),
    .B1(net240),
    .Y(net543));
 sky130_fd_sc_hd__a31oi_1 merge772 (.A1(net129),
    .A2(net861),
    .A3(net44),
    .B1(net232),
    .Y(net544));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(net87),
    .A1(net827),
    .A2(net716),
    .A3(net163),
    .S0(net875),
    .S1(net859),
    .X(net545));
 sky130_fd_sc_hd__mux4_4 merge774 (.A0(net129),
    .A1(net126),
    .A2(net128),
    .A3(net122),
    .S0(net820),
    .S1(net607),
    .X(net546));
 sky130_fd_sc_hd__mux4_1 merge775 (.A0(net216),
    .A1(net213),
    .A2(net202),
    .A3(net214),
    .S0(net218),
    .S1(net912),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 merge776 (.A0(net218),
    .A1(net31),
    .A2(net122),
    .A3(net145),
    .S0(net154),
    .S1(net51),
    .X(net548));
 sky130_fd_sc_hd__mux4_1 merge777 (.A0(net149),
    .A1(net861),
    .A2(net145),
    .A3(net714),
    .S0(net278),
    .S1(net821),
    .X(net549));
 sky130_fd_sc_hd__mux4_4 merge778 (.A0(net437),
    .A1(net441),
    .A2(net350),
    .A3(net336),
    .S0(net344),
    .S1(net659),
    .X(net550));
 sky130_fd_sc_hd__a41oi_1 merge779 (.A1(net732),
    .A2(net858),
    .A3(net725),
    .A4(net147),
    .B1(net958),
    .Y(net551));
 sky130_fd_sc_hd__mux4_4 merge780 (.A0(net443),
    .A1(net426),
    .A2(net349),
    .A3(net120),
    .S0(net338),
    .S1(net658),
    .X(net552));
 sky130_fd_sc_hd__mux4_1 merge781 (.A0(net232),
    .A1(net103),
    .A2(net204),
    .A3(clknet_1_0__leaf_net378),
    .S0(net277),
    .S1(net608),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(net122),
    .A1(net959),
    .A2(net327),
    .A3(net342),
    .S0(net326),
    .S1(net337),
    .X(net554));
 sky130_fd_sc_hd__mux4_4 merge783 (.A0(net341),
    .A1(net335),
    .A2(net337),
    .A3(net244),
    .S0(net242),
    .S1(net115),
    .X(net555));
 sky130_fd_sc_hd__dfrbp_1 merge784 (.CLK(clknet_4_7_0_clk),
    .D(net484),
    .RESET_B(net488),
    .Q(net557),
    .Q_N(net556));
 sky130_fd_sc_hd__dfrbp_2 merge785 (.CLK(clknet_4_2_0_clk),
    .D(net243),
    .RESET_B(net544),
    .Q(net559),
    .Q_N(net558));
 sky130_fd_sc_hd__dfrtn_1 merge786 (.CLK_N(clknet_4_8_0_clk),
    .D(net170),
    .RESET_B(net182),
    .Q(net560));
 sky130_fd_sc_hd__dfrtp_4 merge787 (.CLK(clknet_4_0_0_clk),
    .D(net537),
    .RESET_B(net547),
    .Q(net561));
 sky130_fd_sc_hd__dfrtp_1 merge788 (.CLK(clknet_4_15_0_clk),
    .D(net410),
    .RESET_B(net421),
    .Q(net562));
 sky130_fd_sc_hd__dfrtp_1 merge789 (.CLK(clknet_4_9_0_clk),
    .D(net285),
    .RESET_B(net286),
    .Q(net563));
 sky130_fd_sc_hd__xnor2_1 merge790 (.A(net386),
    .B(net387),
    .Y(net564));
 sky130_fd_sc_hd__xor2_1 merge791 (.A(net370),
    .B(net371),
    .X(net565));
 sky130_fd_sc_hd__dfsbp_2 merge792 (.CLK(clknet_4_2_0_clk),
    .SET_B(net43),
    .Q(net45),
    .Q_N(net566));
 sky130_fd_sc_hd__xnor2_1 merge793 (.A(net297),
    .B(net298),
    .Y(net568));
 sky130_fd_sc_hd__xnor2_1 merge794 (.A(net137),
    .B(net538),
    .Y(net569));
 sky130_fd_sc_hd__xnor2_2 merge795 (.A(net533),
    .B(net522),
    .Y(net570));
 sky130_fd_sc_hd__xor2_1 merge796 (.A(net316),
    .B(net331),
    .X(net571));
 sky130_fd_sc_hd__dfsbp_2 merge797 (.CLK(clknet_4_0_0_clk),
    .SET_B(net118),
    .Q(net573),
    .Q_N(net119));
 sky130_fd_sc_hd__dfstp_1 merge798 (.CLK(clknet_4_10_0_clk),
    .D(net186),
    .SET_B(net192),
    .Q(net828));
 sky130_fd_sc_hd__dfstp_2 merge799 (.CLK(clknet_4_10_0_clk),
    .D(net545),
    .SET_B(net90),
    .Q(net574));
 sky130_fd_sc_hd__xor2_1 merge800 (.A(net64),
    .B(net67),
    .X(net575));
 sky130_fd_sc_hd__dfstp_1 merge801 (.CLK(clknet_4_8_0_clk),
    .D(net157),
    .SET_B(net549),
    .Q(net576));
 sky130_fd_sc_hd__dlrbn_1 merge802 (.D(net515),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net518),
    .Q(net578),
    .Q_N(net577));
 sky130_fd_sc_hd__dlrbn_1 merge803 (.D(net263),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net270),
    .Q(net580),
    .Q_N(net579));
 sky130_fd_sc_hd__dlrbp_2 merge804 (.D(net354),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net534),
    .Q(net582),
    .Q_N(net581));
 sky130_fd_sc_hd__dlrbp_1 merge805 (.D(net449),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net463),
    .Q(net584),
    .Q_N(net583));
 sky130_fd_sc_hd__dlrtn_1 merge806 (.D(net436),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net536),
    .Q(net585));
 sky130_fd_sc_hd__dlrtn_1 merge807 (.D(net380),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net332),
    .Q(net586));
 sky130_fd_sc_hd__xor2_1 merge808 (.A(net469),
    .B(net494),
    .X(net587));
 sky130_fd_sc_hd__dlrtn_1 merge809 (.D(net543),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net546),
    .Q(net588));
 sky130_fd_sc_hd__dlrtp_2 merge810 (.D(net548),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net553),
    .Q(net589));
 sky130_fd_sc_hd__dlrtp_1 merge811 (.D(net400),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net424),
    .Q(net590));
 sky130_fd_sc_hd__dlrtp_2 merge812 (.D(net85),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net66),
    .Q(net835));
 sky130_fd_sc_hd__edfxbp_1 merge813 (.CLK(clknet_4_8_0_clk),
    .D(net575),
    .DE(net68),
    .Q(net592),
    .Q_N(net591));
 sky130_fd_sc_hd__edfxtp_1 merge814 (.CLK(clknet_4_1_0_clk),
    .D(net555),
    .DE(net554),
    .Q(net593));
 sky130_fd_sc_hd__sdlclkp_1 merge815 (.CLK(clknet_4_13_0_clk),
    .GATE(net495),
    .SCE(net532),
    .GCLK(net594));
 sky130_fd_sc_hd__sdlclkp_2 merge816 (.CLK(clknet_4_4_0_clk),
    .GATE(net471),
    .SCE(net550),
    .GCLK(net595));
 sky130_fd_sc_hd__sdlclkp_4 merge817 (.CLK(clknet_4_15_0_clk),
    .GATE(net570),
    .SCE(net528),
    .GCLK(net596));
 sky130_fd_sc_hd__dfrbp_1 merge818 (.CLK(clknet_4_1_0_clk),
    .D(net571),
    .RESET_B(net587),
    .Q(net598),
    .Q_N(net597));
 sky130_fd_sc_hd__xnor2_1 merge819 (.A(net403),
    .B(net422),
    .Y(net599));
 sky130_fd_sc_hd__dfrbp_1 merge820 (.CLK(clknet_4_15_0_clk),
    .D(net299),
    .RESET_B(net527),
    .Q(net601),
    .Q_N(net600));
 sky130_fd_sc_hd__dfrtn_1 merge821 (.CLK_N(clknet_4_11_0_clk),
    .D(net7),
    .RESET_B(net193),
    .Q(net810));
 sky130_fd_sc_hd__dfrtp_4 merge822 (.CLK(clknet_4_11_0_clk),
    .D(net161),
    .RESET_B(net568),
    .Q(net800));
 sky130_fd_sc_hd__dfrtp_1 merge823 (.CLK(clknet_4_15_0_clk),
    .D(net523),
    .RESET_B(net524),
    .Q(net602));
 sky130_fd_sc_hd__dfrtp_1 merge824 (.CLK(clknet_4_6_0_clk),
    .D(net565),
    .RESET_B(net599),
    .Q(net603));
 sky130_fd_sc_hd__dfsbp_1 merge825 (.CLK(clknet_4_8_0_clk),
    .D(net551),
    .SET_B(net166),
    .Q(net605),
    .Q_N(net604));
 sky130_fd_sc_hd__dfsbp_2 merge826 (.CLK(clknet_4_2_0_clk),
    .D(net132),
    .SET_B(net569),
    .Q(net607),
    .Q_N(net606));
 sky130_fd_sc_hd__dfstp_1 merge827 (.CLK(clknet_4_12_0_clk),
    .D(net287),
    .SET_B(net564),
    .Q(net608));
 sky130_fd_sc_hd__dfstp_1 merge828 (.CLK(clknet_4_10_0_clk),
    .D(net97),
    .Q(net845));
 sky130_fd_sc_hd__dfxbp_1 s829 (.CLK(clknet_4_10_0_clk),
    .D(net160),
    .Q(net610),
    .Q_N(net609));
 sky130_fd_sc_hd__dfxbp_1 s830 (.CLK(clknet_4_10_0_clk),
    .D(net171),
    .Q(net612),
    .Q_N(net611));
 sky130_fd_sc_hd__dfxtp_1 s831 (.CLK(clknet_4_9_0_clk),
    .D(net181),
    .Q(net613));
 sky130_fd_sc_hd__dfxtp_2 s832 (.CLK(clknet_4_10_0_clk),
    .D(net183),
    .Q(net614));
 sky130_fd_sc_hd__dfxtp_2 s833 (.CLK(clknet_4_10_0_clk),
    .D(net187),
    .Q(net615));
 sky130_fd_sc_hd__dlclkp_1 s834 (.CLK(clknet_4_11_0_clk),
    .GATE(net188),
    .GCLK(net616));
 sky130_fd_sc_hd__dlclkp_2 s835 (.CLK(clknet_4_10_0_clk),
    .GATE(net194),
    .GCLK(net617));
 sky130_fd_sc_hd__dlclkp_4 s836 (.CLK(clknet_4_11_0_clk),
    .GATE(net195),
    .GCLK(net803));
 sky130_fd_sc_hd__dlxbn_1 s837 (.D(net198),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net819),
    .Q_N(net618));
 sky130_fd_sc_hd__dlxbn_1 s838 (.D(net199),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net620),
    .Q_N(net619));
 sky130_fd_sc_hd__dlxbp_1 s839 (.D(net219),
    .GATE(clknet_4_0_0_clk),
    .Q(net622),
    .Q_N(net621));
 sky130_fd_sc_hd__dlxtn_4 s840 (.D(net222),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net623));
 sky130_fd_sc_hd__dlxtn_2 s841 (.D(net241),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net624));
 sky130_fd_sc_hd__dlxtn_1 s842 (.D(net295),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net625));
 sky130_fd_sc_hd__dlxtp_1 s843 (.D(net301),
    .GATE(clknet_4_14_0_clk),
    .Q(net626));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s844 (.D(net302),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net627));
 sky130_fd_sc_hd__dfxbp_1 s845 (.CLK(clknet_4_14_0_clk),
    .D(net308),
    .Q(net629),
    .Q_N(net628));
 sky130_fd_sc_hd__dfxbp_1 s846 (.CLK(clknet_4_12_0_clk),
    .D(net328),
    .Q(net631),
    .Q_N(net630));
 sky130_fd_sc_hd__dfxtp_1 s847 (.CLK(clknet_4_1_0_clk),
    .D(net330),
    .Q(net632));
 sky130_fd_sc_hd__dfxtp_2 s848 (.CLK(clknet_4_6_0_clk),
    .D(net345),
    .Q(net633));
 sky130_fd_sc_hd__dfxtp_2 s849 (.CLK(clknet_4_6_0_clk),
    .D(net356),
    .Q(net634));
 sky130_fd_sc_hd__dlclkp_1 s850 (.CLK(clknet_4_6_0_clk),
    .GATE(net372),
    .GCLK(net635));
 sky130_fd_sc_hd__dlclkp_2 s851 (.CLK(clknet_4_3_0_clk),
    .GATE(net373),
    .GCLK(net636));
 sky130_fd_sc_hd__dlclkp_4 s852 (.CLK(clknet_4_3_0_clk),
    .GATE(net374),
    .GCLK(net637));
 sky130_fd_sc_hd__dlxbn_1 s853 (.D(net376),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net639),
    .Q_N(net638));
 sky130_fd_sc_hd__dlxbn_2 s854 (.D(net381),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net641),
    .Q_N(net640));
 sky130_fd_sc_hd__dlxbp_1 s855 (.D(net382),
    .GATE(clknet_4_6_0_clk),
    .Q(net643),
    .Q_N(net642));
 sky130_fd_sc_hd__dlxtn_1 s856 (.D(net398),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net791));
 sky130_fd_sc_hd__dlxtn_2 s857 (.D(net401),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net644));
 sky130_fd_sc_hd__dlxtn_2 s858 (.D(net402),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net645));
 sky130_fd_sc_hd__dlxtp_1 s859 (.D(net405),
    .GATE(clknet_4_13_0_clk),
    .Q(net646));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s860 (.D(net407),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net647));
 sky130_fd_sc_hd__dfxbp_1 s861 (.CLK(clknet_4_14_0_clk),
    .D(net408),
    .Q(net649),
    .Q_N(net648));
 sky130_fd_sc_hd__dfxbp_1 s862 (.CLK(clknet_4_14_0_clk),
    .D(net411),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__dfxtp_1 s863 (.CLK(clknet_4_12_0_clk),
    .D(net412),
    .Q(net652));
 sky130_fd_sc_hd__dfxtp_2 s864 (.CLK(clknet_4_14_0_clk),
    .D(net413),
    .Q(net653));
 sky130_fd_sc_hd__dfxtp_2 s865 (.CLK(clknet_4_15_0_clk),
    .D(net415),
    .Q(net654));
 sky130_fd_sc_hd__dlclkp_1 s866 (.CLK(clknet_4_14_0_clk),
    .GATE(net416),
    .GCLK(net655));
 sky130_fd_sc_hd__dlclkp_2 s867 (.CLK(clknet_4_15_0_clk),
    .GATE(net420),
    .GCLK(net656));
 sky130_fd_sc_hd__dlclkp_4 s868 (.CLK(clknet_4_13_0_clk),
    .GATE(net425),
    .GCLK(net657));
 sky130_fd_sc_hd__dlxbn_1 s869 (.D(net440),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net659),
    .Q_N(net658));
 sky130_fd_sc_hd__dlxbn_2 s870 (.D(net446),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net661),
    .Q_N(net660));
 sky130_fd_sc_hd__dlxbp_1 s871 (.D(net466),
    .GATE(clknet_4_5_0_clk),
    .Q(net663),
    .Q_N(net662));
 sky130_fd_sc_hd__dlxtn_2 s872 (.D(net468),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net664));
 sky130_fd_sc_hd__dlxtn_1 s873 (.D(net470),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net665));
 sky130_fd_sc_hd__dlxtn_1 s874 (.D(net475),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net666));
 sky130_fd_sc_hd__dlxtp_1 s875 (.D(net481),
    .GATE(clknet_4_7_0_clk),
    .Q(net667));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s876 (.D(net482),
    .SLEEP_B(clknet_4_7_0_clk),
    .Q(net668));
 sky130_fd_sc_hd__dfxbp_1 s877 (.CLK(clknet_4_7_0_clk),
    .D(net485),
    .Q(net670),
    .Q_N(net669));
 sky130_fd_sc_hd__dfxbp_1 s878 (.CLK(clknet_4_7_0_clk),
    .D(net490),
    .Q(net672),
    .Q_N(net671));
 sky130_fd_sc_hd__dfxtp_1 s879 (.CLK(clknet_4_7_0_clk),
    .D(net491),
    .Q(net673));
 sky130_fd_sc_hd__dfxtp_1 s880 (.CLK(clknet_4_7_0_clk),
    .D(net492),
    .Q(net674));
 sky130_fd_sc_hd__dfxtp_1 s881 (.CLK(clknet_4_13_0_clk),
    .D(net503),
    .Q(net675));
 sky130_fd_sc_hd__dlclkp_1 s882 (.CLK(clknet_4_13_0_clk),
    .GATE(net509),
    .GCLK(net676));
 sky130_fd_sc_hd__dlclkp_2 s883 (.CLK(clknet_4_13_0_clk),
    .GATE(net520),
    .GCLK(net677));
 sky130_fd_sc_hd__dlclkp_4 s884 (.CLK(clknet_4_15_0_clk),
    .GATE(net530),
    .GCLK(net678));
 sky130_fd_sc_hd__dlxbn_1 s885 (.D(net535),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net680),
    .Q_N(net679));
 sky130_fd_sc_hd__dlxbn_1 s886 (.D(net542),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dlxbp_1 s887 (.D(net552),
    .GATE(clknet_4_4_0_clk),
    .Q(net684),
    .Q_N(net683));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(in0),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net685));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net686));
 sky130_fd_sc_hd__buf_1 input4 (.A(in11),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(in12),
    .X(net688));
 sky130_fd_sc_hd__buf_12 input6 (.A(in13),
    .X(net689));
 sky130_fd_sc_hd__buf_4 input7 (.A(in14),
    .X(net690));
 sky130_fd_sc_hd__buf_1 input8 (.A(in15),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_8 input9 (.A(in16),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net693));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(in18),
    .X(net694));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(in19),
    .X(net695));
 sky130_fd_sc_hd__buf_2 input13 (.A(in2),
    .X(net696));
 sky130_fd_sc_hd__buf_1 input14 (.A(in20),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(in21),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(in22),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(in23),
    .X(net700));
 sky130_fd_sc_hd__buf_4 input18 (.A(in24),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in25),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_8 input20 (.A(in26),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(in27),
    .X(net704));
 sky130_fd_sc_hd__buf_2 input22 (.A(in28),
    .X(net705));
 sky130_fd_sc_hd__buf_4 input23 (.A(in29),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(in3),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_8 input26 (.A(in31),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(in33),
    .X(net711));
 sky130_fd_sc_hd__buf_1 input29 (.A(in34),
    .X(net712));
 sky130_fd_sc_hd__buf_1 input30 (.A(in35),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(in36),
    .X(net714));
 sky130_fd_sc_hd__buf_1 input32 (.A(in37),
    .X(net715));
 sky130_fd_sc_hd__buf_4 input33 (.A(in38),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(in39),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_8 input35 (.A(in4),
    .X(net718));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net719));
 sky130_fd_sc_hd__buf_1 input37 (.A(in41),
    .X(net720));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(in43),
    .X(net722));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(in44),
    .X(net723));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net724));
 sky130_fd_sc_hd__buf_4 input42 (.A(in46),
    .X(net725));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(in47),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net727));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(in5),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(in50),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in51),
    .X(net731));
 sky130_fd_sc_hd__buf_1 input49 (.A(in52),
    .X(net732));
 sky130_fd_sc_hd__buf_1 input50 (.A(in53),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net734));
 sky130_fd_sc_hd__buf_1 input52 (.A(in55),
    .X(net735));
 sky130_fd_sc_hd__buf_2 input53 (.A(in56),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in57),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(in58),
    .X(net738));
 sky130_fd_sc_hd__buf_1 input56 (.A(in6),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(in60),
    .X(net740));
 sky130_fd_sc_hd__buf_1 input58 (.A(in61),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(in62),
    .X(net742));
 sky130_fd_sc_hd__buf_1 input60 (.A(in63),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(in64),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(in65),
    .X(net745));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(in66),
    .X(net746));
 sky130_fd_sc_hd__buf_1 input64 (.A(in67),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(in68),
    .X(net748));
 sky130_fd_sc_hd__buf_1 input66 (.A(in69),
    .X(net749));
 sky130_fd_sc_hd__buf_4 input67 (.A(in7),
    .X(net750));
 sky130_fd_sc_hd__buf_1 input68 (.A(in70),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(in71),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(in72),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(in73),
    .X(net754));
 sky130_fd_sc_hd__buf_1 input72 (.A(in74),
    .X(net755));
 sky130_fd_sc_hd__buf_1 input73 (.A(in75),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(in76),
    .X(net757));
 sky130_fd_sc_hd__buf_1 input75 (.A(in77),
    .X(net758));
 sky130_fd_sc_hd__buf_1 input76 (.A(in78),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(in79),
    .X(net760));
 sky130_fd_sc_hd__buf_4 input78 (.A(in8),
    .X(net761));
 sky130_fd_sc_hd__buf_1 input79 (.A(in80),
    .X(net762));
 sky130_fd_sc_hd__dlymetal6s2s_1 input80 (.A(in81),
    .X(net763));
 sky130_fd_sc_hd__buf_1 input81 (.A(in82),
    .X(net764));
 sky130_fd_sc_hd__dlymetal6s2s_1 input82 (.A(in83),
    .X(net765));
 sky130_fd_sc_hd__buf_1 input83 (.A(in84),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(in85),
    .X(net767));
 sky130_fd_sc_hd__buf_1 input85 (.A(in86),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(in87),
    .X(net769));
 sky130_fd_sc_hd__buf_1 input87 (.A(in88),
    .X(net770));
 sky130_fd_sc_hd__buf_1 input88 (.A(in89),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(in9),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(in90),
    .X(net773));
 sky130_fd_sc_hd__buf_2 input91 (.A(in91),
    .X(net774));
 sky130_fd_sc_hd__buf_1 input92 (.A(in92),
    .X(net775));
 sky130_fd_sc_hd__buf_1 input93 (.A(in93),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_4 input94 (.A(in94),
    .X(net777));
 sky130_fd_sc_hd__buf_4 input95 (.A(in95),
    .X(net778));
 sky130_fd_sc_hd__buf_2 input96 (.A(in96),
    .X(net779));
 sky130_fd_sc_hd__buf_1 input97 (.A(in97),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(in98),
    .X(net781));
 sky130_fd_sc_hd__buf_1 input99 (.A(in99),
    .X(net782));
 sky130_fd_sc_hd__buf_2 output100 (.A(net783),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net784),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net785),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net786),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net787),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output105 (.A(net788),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net789),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output107 (.A(net790),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output108 (.A(net791),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net792),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net793),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output111 (.A(net794),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output112 (.A(net859),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net796),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net797),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(clknet_1_1__leaf_net798),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net799),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net800),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net801),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net802),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(clknet_1_1__leaf_net803),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output121 (.A(net804),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_4 output122 (.A(net805),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_4 output123 (.A(net806),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(clknet_1_1__leaf_net807),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net442),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net809),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net810),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net811),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net812),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_4 output130 (.A(net813),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output131 (.A(net874),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output132 (.A(net815),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net816),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_4 output134 (.A(net817),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_4 output135 (.A(net818),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_4 output136 (.A(net819),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output137 (.A(net820),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output138 (.A(net821),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(clknet_1_1__leaf_net822),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net823),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net824),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output142 (.A(net825),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net826),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output144 (.A(net827),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net828),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_4 output146 (.A(net829),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output147 (.A(net830),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_4 output148 (.A(net831),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output149 (.A(net832),
    .X(out63));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net833),
    .X(out64));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(clknet_1_1__leaf_net834),
    .X(out65));
 sky130_fd_sc_hd__buf_2 output152 (.A(net835),
    .X(out69));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net836),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net837),
    .X(out73));
 sky130_fd_sc_hd__clkbuf_4 output155 (.A(net838),
    .X(out75));
 sky130_fd_sc_hd__buf_2 output156 (.A(net839),
    .X(out78));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(clknet_1_1__leaf_net840),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output158 (.A(net841),
    .X(out80));
 sky130_fd_sc_hd__clkbuf_4 output159 (.A(net842),
    .X(out81));
 sky130_fd_sc_hd__buf_2 output160 (.A(net843),
    .X(out84));
 sky130_fd_sc_hd__buf_2 output161 (.A(net844),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output162 (.A(net845),
    .X(out87));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net846),
    .X(out88));
 sky130_fd_sc_hd__clkbuf_4 output164 (.A(net847),
    .X(out89));
 sky130_fd_sc_hd__clkbuf_4 output165 (.A(net848),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 output166 (.A(net849),
    .X(out90));
 sky130_fd_sc_hd__clkbuf_4 output167 (.A(net850),
    .X(out91));
 sky130_fd_sc_hd__clkbuf_4 output168 (.A(net851),
    .X(out92));
 sky130_fd_sc_hd__clkbuf_4 output169 (.A(net852),
    .X(out93));
 sky130_fd_sc_hd__clkbuf_4 output170 (.A(net853),
    .X(out95));
 sky130_fd_sc_hd__clkbuf_4 output171 (.A(net854),
    .X(out96));
 sky130_fd_sc_hd__clkbuf_4 output172 (.A(net855),
    .X(out97));
 sky130_fd_sc_hd__buf_8 fanout173 (.A(net817),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_4 fanout174 (.A(net432),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_4 max_cap175 (.A(net63),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_8 fanout176 (.A(net795),
    .X(net859));
 sky130_fd_sc_hd__buf_4 fanout177 (.A(net429),
    .X(net860));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net41),
    .X(net861));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net426),
    .X(net862));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(net315),
    .X(net863));
 sky130_fd_sc_hd__buf_2 max_cap181 (.A(net58),
    .X(net864));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(net786),
    .X(net865));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(net841),
    .X(net866));
 sky130_fd_sc_hd__buf_4 max_cap184 (.A(net28),
    .X(net867));
 sky130_fd_sc_hd__buf_4 max_cap185 (.A(net208),
    .X(net868));
 sky130_fd_sc_hd__buf_4 max_cap186 (.A(net788),
    .X(net869));
 sky130_fd_sc_hd__buf_8 fanout187 (.A(net56),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_4 max_cap188 (.A(net25),
    .X(net871));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net53),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net53),
    .X(net873));
 sky130_fd_sc_hd__buf_8 fanout191 (.A(net814),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net876),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(net877),
    .X(net876));
 sky130_fd_sc_hd__buf_2 fanout194 (.A(net879),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(net879),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_4 fanout196 (.A(net167),
    .X(net879));
 sky130_fd_sc_hd__buf_4 max_cap197 (.A(net19),
    .X(net880));
 sky130_fd_sc_hd__buf_4 max_cap198 (.A(net17),
    .X(net881));
 sky130_fd_sc_hd__clkbuf_4 fanout199 (.A(net156),
    .X(net882));
 sky130_fd_sc_hd__buf_4 max_cap200 (.A(net12),
    .X(net883));
 sky130_fd_sc_hd__buf_12 wire201 (.A(net8),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(net667),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_4 fanout203 (.A(net770),
    .X(net886));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(net765),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(net765),
    .X(net888));
 sky130_fd_sc_hd__buf_4 fanout206 (.A(net763),
    .X(net889));
 sky130_fd_sc_hd__buf_12 fanout207 (.A(net892),
    .X(net890));
 sky130_fd_sc_hd__buf_2 fanout208 (.A(net892),
    .X(net891));
 sky130_fd_sc_hd__buf_12 fanout209 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__buf_12 fanout210 (.A(net689),
    .X(net893));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_4 fanout212 (.A(net733),
    .X(net895));
 sky130_fd_sc_hd__buf_2 max_cap213 (.A(net283),
    .X(net896));
 sky130_fd_sc_hd__inv_16 c676_1 (.A(clknet_1_1__leaf_net595),
    .Y(net897));
 sky130_fd_sc_hd__inv_16 net799_2 (.A(clknet_1_1__leaf_net595),
    .Y(net898));
 sky130_fd_sc_hd__inv_16 net898_3 (.A(clknet_1_1__leaf_net595),
    .Y(net899));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net678 (.A(net678),
    .X(clknet_0_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net678 (.A(clknet_0_net678),
    .X(clknet_1_0__leaf_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net678 (.A(clknet_0_net678),
    .X(clknet_1_1__leaf_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net596 (.A(net596),
    .X(clknet_0_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_1__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net594 (.A(net594),
    .X(clknet_0_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net594 (.A(clknet_0_net594),
    .X(clknet_1_0__leaf_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net594 (.A(clknet_0_net594),
    .X(clknet_1_1__leaf_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net496 (.A(net496),
    .X(clknet_0_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_0__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_1__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net505 (.A(net505),
    .X(clknet_0_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net505 (.A(clknet_0_net505),
    .X(clknet_1_0__leaf_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net505 (.A(clknet_0_net505),
    .X(clknet_1_1__leaf_net505));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net517 (.A(net517),
    .X(clknet_0_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_0__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_1__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net499 (.A(net499),
    .X(clknet_0_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_0__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_1__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net676 (.A(net676),
    .X(clknet_0_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_0__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_1__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net677 (.A(net677),
    .X(clknet_0_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_0__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_1__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net526 (.A(net526),
    .X(clknet_0_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_0__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_1__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net521 (.A(net521),
    .X(clknet_0_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_0__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_1__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net497 (.A(net497),
    .X(clknet_0_net497));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net497 (.A(clknet_0_net497),
    .X(clknet_1_0__leaf_net497));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net497 (.A(clknet_0_net497),
    .X(clknet_1_1__leaf_net497));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net504 (.A(net504),
    .X(clknet_0_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_0__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_1__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net513 (.A(net513),
    .X(clknet_0_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_0__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_1__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net657 (.A(net657),
    .X(clknet_0_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_0__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_1__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net656 (.A(net656),
    .X(clknet_0_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_0__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_1__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net423 (.A(net423),
    .X(clknet_0_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_0__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_1__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net655 (.A(net655),
    .X(clknet_0_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net418 (.A(net418),
    .X(clknet_0_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net418 (.A(clknet_0_net418),
    .X(clknet_1_0__leaf_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net418 (.A(clknet_0_net418),
    .X(clknet_1_1__leaf_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net637 (.A(net637),
    .X(clknet_0_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net637 (.A(clknet_0_net637),
    .X(clknet_1_0__leaf_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net637 (.A(clknet_0_net637),
    .X(clknet_1_1__leaf_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net404 (.A(net404),
    .X(clknet_0_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net393 (.A(net393),
    .X(clknet_0_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net393 (.A(clknet_0_net393),
    .X(clknet_1_0__leaf_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net393 (.A(clknet_0_net393),
    .X(clknet_1_1__leaf_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net377 (.A(net377),
    .X(clknet_0_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_0__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_1__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net378 (.A(net378),
    .X(clknet_0_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_1__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net636 (.A(net636),
    .X(clknet_0_net636));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net636 (.A(clknet_0_net636),
    .X(clknet_1_0__leaf_net636));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net636 (.A(clknet_0_net636),
    .X(clknet_1_1__leaf_net636));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net635 (.A(net635),
    .X(clknet_0_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net635 (.A(clknet_0_net635),
    .X(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net635 (.A(clknet_0_net635),
    .X(clknet_1_1__leaf_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net803 (.A(net803),
    .X(clknet_0_net803));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net803 (.A(clknet_0_net803),
    .X(clknet_1_0__leaf_net803));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net803 (.A(clknet_0_net803),
    .X(clknet_1_1__leaf_net803));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net617 (.A(net617),
    .X(clknet_0_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net617 (.A(clknet_0_net617),
    .X(clknet_1_0__leaf_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net617 (.A(clknet_0_net617),
    .X(clknet_1_1__leaf_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net807 (.A(net807),
    .X(clknet_0_net807));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net807 (.A(clknet_0_net807),
    .X(clknet_1_0__leaf_net807));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net807 (.A(clknet_0_net807),
    .X(clknet_1_1__leaf_net807));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net798 (.A(net798),
    .X(clknet_0_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_0__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_1__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net616 (.A(net616),
    .X(clknet_0_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_0__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_1__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net834 (.A(net834),
    .X(clknet_0_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_0__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net822 (.A(net822),
    .X(clknet_0_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net822 (.A(clknet_0_net822),
    .X(clknet_1_0__leaf_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net822 (.A(net905),
    .X(clknet_1_1__leaf_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net200 (.A(net200),
    .X(clknet_0_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_0__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net200 (.A(net907),
    .X(clknet_1_1__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net840 (.A(net840),
    .X(clknet_0_net840));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net840 (.A(clknet_0_net840),
    .X(clknet_1_0__leaf_net840));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net840 (.A(clknet_0_net840),
    .X(clknet_1_1__leaf_net840));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net309 (.A(net309),
    .X(clknet_0_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net309 (.A(clknet_0_net309),
    .X(clknet_1_0__leaf_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net309 (.A(clknet_0_net309),
    .X(clknet_1_1__leaf_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net303 (.A(net303),
    .X(clknet_0_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_0__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net303 (.A(clknet_0_net303),
    .X(clknet_1_1__leaf_net303));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net189 (.A(net189),
    .X(clknet_0_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_0__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net189 (.A(clknet_0_net189),
    .X(clknet_1_1__leaf_net189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net483 (.A(net483),
    .X(clknet_0_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net483 (.A(clknet_0_net483),
    .X(clknet_1_0__leaf_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net483 (.A(clknet_0_net483),
    .X(clknet_1_1__leaf_net483));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net472 (.A(net472),
    .X(clknet_0_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_0__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net472 (.A(clknet_0_net472),
    .X(clknet_1_1__leaf_net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net355 (.A(net355),
    .X(clknet_0_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_0__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_1__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net808),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net845),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net59),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net82),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_1 clone5 (.A(net56),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer6 (.A(net56),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(clknet_0_net822),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_1 clone8 (.A(net892),
    .X(net906));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer9 (.A(clknet_0_net200),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_1 clone10 (.A(net817),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net825),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net909),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net433),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net621),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net663),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net174),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net634),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net614),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net835),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net579),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net632),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net580),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net576),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net793),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net133),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net625),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net320),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net293),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net612),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net683),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net224),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net253),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net250),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net668),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net563),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net258),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net126),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net613),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net322),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net633),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net643),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net672),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net660),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net305),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net333),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net674),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net294),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net674),
    .X(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B1_N (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_RESET_B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_Y (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A4 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B1_N (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_SCE (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_Y (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B1_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_Y (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_S1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B1_N (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A4 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_SET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_D (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_Y (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A3 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_SCD (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_Y (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_D (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B1_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B1_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_D (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Y (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_SCE (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_SCD (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_SCE (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_Q (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCE (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_SCE (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_Q_N (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B1_N (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A0 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A0 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A4 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_SCE (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B1_N (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_Q_N (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A4 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_X (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_Y (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_D (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B1_N (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_SCD (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_Y (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A0 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_RESET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_X (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_X (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap197_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_Y (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A4 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SCE (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_Y (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_D (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_SCE (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A3 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B1_N (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B1_N (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_Y (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_B1_N (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_S1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_Y (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A3 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_SCD (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A3 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_S0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_Y (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_Y (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_SCE (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_D (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_X (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_RESET_B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_SCE (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_SCD (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_X (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_Y (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A0 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SET_B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_Q (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_Q_N (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_S0 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_Q_N (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_SCD (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_X (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_Q (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_Y (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_D (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_Y (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_D (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_Y (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_RESET_B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S0 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A0 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_Y (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_Y (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A3 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_SCE (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_Y (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold39_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A4 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_Q_N (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_Q (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_DE (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_SCD (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_Y (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_SCD (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_SET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_SCD (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_Y (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_s846_D (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_X (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A3 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_Y (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_S1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_Y (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B1_N (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_Y (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_SCE (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCD (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_Y (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A3 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_Y (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_SCE (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_X (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_SCE (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A4 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_Q_N (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_Q (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_D (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_X (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_DE (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_X (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_SCD (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_X (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_X (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_B1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_RESET_B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_Q (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCE (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_Q_N (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_Q (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_X (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_Q_N (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_SCE (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1_N (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B1_N (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_Q (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_Q (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A3 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_Q_N (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A4 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_Q (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_S1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SCE (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_s829_Q (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_SCE (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_B1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold18_A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_s832_Q (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_SET_B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_s838_Q_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_s838_Q (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_s840_Q (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_SCE (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCE (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1_N (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_SET_B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_Q (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_B1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_B1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_B1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_Q_N (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_Q (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_Q (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_Q_N (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_Q (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_Q (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_Q (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B1_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_SCE (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_B1_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_D (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_SCD (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire201_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SCD (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_Y (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A3 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A3 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_X (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_RESET_B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_Y (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_S (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B1_N (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A2 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1_N (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A0 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_SCE (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A3 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_SCD (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_S0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A4 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A3 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A4 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_RESET_B (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A2 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B1_N (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A3 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_SCD (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1_N (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A2 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B1_N (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A4 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S0 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B1_N (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A3 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_S1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A4 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_X (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S0 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_B1_N (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A0 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A3 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A0 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A4 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_X (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_X (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A3 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A2 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A3 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_X (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCD (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_SCE (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A2 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_Q (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_Q (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_X (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A4 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap186_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_Y (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B1_N (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Y (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A4 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_Q (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold24_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_Q (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_SCD (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_SCD (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_Q (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B1_N (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_RESET_B (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_Y (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A4 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_RESET_B (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_Q (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_Q (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_Y (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_SET_B (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_SCE (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_SCD (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_Y (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_S1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_B1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_Y (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_Y (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_Y (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_Y (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A4 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A4 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_Y (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_B1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_SCE (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SET_B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A4 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A3 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_S0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap175_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCD (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_SCE (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A4 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_SET_B (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SCD (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_RESET_B (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_B1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_SCD (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_SCE (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A4 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A4 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_RESET_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B1_N (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_SCD (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A4 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_SET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap181_X (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B1_N (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_SCD (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_RESET_B (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_SET_B (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap184_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap185_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap186_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_SCD (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A2 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap188_X (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A4 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B1_N (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A4 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A4 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A4 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A4 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A4 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A4 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_SCE (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap197_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap198_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_SCE (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap200_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_S1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire201_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_SCE (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B1_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_RESET_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A4 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_SCD (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B1_N (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B1_N (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_S (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B1_N (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_SET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone8_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_B1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_SET_B (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCE (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_SCE (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s839_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s840_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s831_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s834_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s836_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s837_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s838_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s842_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s846_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A4 (.DIODE(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A3 (.DIODE(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net378_X (.DIODE(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone5_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_SCD (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_RESET_B (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_RESET_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_SET_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold37_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net125));
 sky130_fd_sc_hd__clkbuf_1 clone1 (.A(net8),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net20),
    .X(net948));
 sky130_fd_sc_hd__a31o_1 clone6 (.A1(net96),
    .A2(net92),
    .A3(net592),
    .B1(net845),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net52),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net950),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net951),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_1 clone14 (.A(net56),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_1 clone15 (.A(net959),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net74),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_1 clone17 (.A(net689),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_1 clone18 (.A(net958),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_1 clone19 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_1 clone20 (.A(net689),
    .X(net959));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
