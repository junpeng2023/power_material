module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire clknet_0_clk;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net714;
 wire clknet_1_0__leaf_net714;
 wire clknet_1_1__leaf_net714;
 wire clknet_0_net360;
 wire clknet_1_0__leaf_net360;
 wire clknet_1_1__leaf_net360;
 wire clknet_0_net410;
 wire clknet_1_0__leaf_net410;
 wire clknet_1_1__leaf_net410;
 wire clknet_0_net404;
 wire clknet_1_0__leaf_net404;
 wire clknet_1_1__leaf_net404;
 wire clknet_0_net378;
 wire clknet_1_0__leaf_net378;
 wire clknet_1_1__leaf_net378;
 wire clknet_0_net417;
 wire clknet_1_0__leaf_net417;
 wire clknet_1_1__leaf_net417;
 wire clknet_0_net627;
 wire clknet_1_0__leaf_net627;
 wire clknet_1_1__leaf_net627;
 wire clknet_0_net333;
 wire clknet_1_0__leaf_net333;
 wire clknet_1_1__leaf_net333;
 wire clknet_0_net355;
 wire clknet_1_0__leaf_net355;
 wire clknet_1_1__leaf_net355;
 wire clknet_0_net477;
 wire clknet_1_0__leaf_net477;
 wire clknet_1_1__leaf_net477;
 wire clknet_0_net361;
 wire clknet_1_0__leaf_net361;
 wire clknet_1_1__leaf_net361;
 wire clknet_0_net368;
 wire clknet_1_0__leaf_net368;
 wire clknet_1_1__leaf_net368;
 wire clknet_0_net694;
 wire clknet_1_0__leaf_net694;
 wire clknet_1_1__leaf_net694;
 wire clknet_0_net381;
 wire clknet_1_0__leaf_net381;
 wire clknet_1_1__leaf_net381;
 wire clknet_0_net858;
 wire clknet_1_0__leaf_net858;
 wire clknet_1_1__leaf_net858;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net371;
 wire clknet_1_0__leaf_net371;
 wire clknet_1_1__leaf_net371;
 wire clknet_0_net369;
 wire clknet_1_0__leaf_net369;
 wire clknet_1_1__leaf_net369;
 wire clknet_0_net359;
 wire clknet_1_0__leaf_net359;
 wire clknet_1_1__leaf_net359;
 wire clknet_0_net382;
 wire clknet_1_0__leaf_net382;
 wire clknet_1_1__leaf_net382;
 wire clknet_0_net383;
 wire clknet_1_0__leaf_net383;
 wire clknet_1_1__leaf_net383;
 wire clknet_0_net695;
 wire clknet_1_0__leaf_net695;
 wire clknet_1_1__leaf_net695;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire clknet_0_net395;
 wire clknet_1_0__leaf_net395;
 wire clknet_1_1__leaf_net395;
 wire clknet_0_net832;
 wire clknet_1_0__leaf_net832;
 wire clknet_1_1__leaf_net832;
 wire clknet_0_net815;
 wire clknet_1_0__leaf_net815;
 wire clknet_1_1__leaf_net815;
 wire clknet_0_net435;
 wire clknet_1_0__leaf_net435;
 wire clknet_1_1__leaf_net435;
 wire clknet_0_net693;
 wire clknet_1_0__leaf_net693;
 wire clknet_1_1__leaf_net693;
 wire clknet_0_net484;
 wire clknet_1_0__leaf_net484;
 wire clknet_1_1__leaf_net484;
 wire clknet_0_net365;
 wire clknet_1_0__leaf_net365;
 wire clknet_1_1__leaf_net365;
 wire clknet_0_net713;
 wire clknet_1_0__leaf_net713;
 wire clknet_1_1__leaf_net713;
 wire clknet_0_net821;
 wire clknet_1_0__leaf_net821;
 wire clknet_1_1__leaf_net821;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire clknet_0_net712;
 wire clknet_1_0__leaf_net712;
 wire clknet_1_1__leaf_net712;
 wire clknet_0_net678;
 wire clknet_1_0__leaf_net678;
 wire clknet_1_1__leaf_net678;
 wire clknet_0_net305;
 wire clknet_1_0__leaf_net305;
 wire clknet_1_1__leaf_net305;
 wire clknet_0_net677;
 wire clknet_1_0__leaf_net677;
 wire clknet_1_1__leaf_net677;
 wire clknet_0_net676;
 wire clknet_1_0__leaf_net676;
 wire clknet_1_1__leaf_net676;
 wire clknet_0_net302;
 wire clknet_1_0__leaf_net302;
 wire clknet_1_1__leaf_net302;
 wire clknet_0_net307;
 wire clknet_1_0__leaf_net307;
 wire clknet_1_1__leaf_net307;
 wire clknet_0_net296;
 wire clknet_1_0__leaf_net296;
 wire clknet_1_1__leaf_net296;
 wire clknet_0_net298;
 wire clknet_1_0__leaf_net298;
 wire clknet_1_1__leaf_net298;
 wire clknet_0_net659;
 wire clknet_1_0__leaf_net659;
 wire clknet_1_1__leaf_net659;
 wire clknet_0_net202;
 wire clknet_1_0__leaf_net202;
 wire clknet_1_1__leaf_net202;
 wire clknet_0_net182;
 wire clknet_1_0__leaf_net182;
 wire clknet_1_1__leaf_net182;
 wire clknet_0_net425;
 wire clknet_1_0__leaf_net425;
 wire clknet_1_1__leaf_net425;
 wire clknet_0_net424;
 wire clknet_1_0__leaf_net424;
 wire clknet_1_1__leaf_net424;
 wire clknet_0_net314;
 wire clknet_1_0__leaf_net314;
 wire clknet_1_1__leaf_net314;
 wire clknet_0_net317;
 wire clknet_1_0__leaf_net317;
 wire clknet_1_1__leaf_net317;
 wire clknet_0_net287;
 wire clknet_1_0__leaf_net287;
 wire clknet_1_1__leaf_net287;
 wire clknet_0_net294;
 wire clknet_1_0__leaf_net294;
 wire clknet_1_1__leaf_net294;
 wire clknet_0_net206;
 wire clknet_1_0__leaf_net206;
 wire clknet_1_1__leaf_net206;
 wire clknet_0_net195;
 wire clknet_1_0__leaf_net195;
 wire clknet_1_1__leaf_net195;
 wire clknet_0_net316;
 wire clknet_1_0__leaf_net316;
 wire clknet_1_1__leaf_net316;
 wire clknet_0_net192;
 wire clknet_1_0__leaf_net192;
 wire clknet_1_1__leaf_net192;
 wire clknet_0_net844;
 wire clknet_1_0__leaf_net844;
 wire clknet_1_1__leaf_net844;
 wire clknet_0_net184;
 wire clknet_1_0__leaf_net184;
 wire clknet_1_1__leaf_net184;
 wire clknet_0_net288;
 wire clknet_1_0__leaf_net288;
 wire clknet_1_1__leaf_net288;
 wire clknet_0_net285;
 wire clknet_1_0__leaf_net285;
 wire clknet_1_1__leaf_net285;
 wire clknet_0_net286;
 wire clknet_1_0__leaf_net286;
 wire clknet_1_1__leaf_net286;
 wire clknet_0_net183;
 wire clknet_1_0__leaf_net183;
 wire clknet_1_1__leaf_net183;
 wire clknet_0_net165;
 wire clknet_1_0__leaf_net165;
 wire clknet_1_1__leaf_net165;
 wire clknet_0_net167;
 wire clknet_1_0__leaf_net167;
 wire clknet_1_1__leaf_net167;
 wire clknet_0_net625;
 wire clknet_1_0__leaf_net625;
 wire clknet_1_1__leaf_net625;
 wire clknet_0_net151;
 wire clknet_1_0__leaf_net151;
 wire clknet_1_1__leaf_net151;
 wire clknet_0_net150;
 wire clknet_1_0__leaf_net150;
 wire clknet_1_1__leaf_net150;
 wire clknet_0_net156;
 wire clknet_1_0__leaf_net156;
 wire clknet_1_1__leaf_net156;
 wire clknet_0_net154;
 wire clknet_1_0__leaf_net154;
 wire clknet_1_1__leaf_net154;
 wire clknet_0_net161;
 wire clknet_1_0__leaf_net161;
 wire clknet_1_1__leaf_net161;
 wire clknet_0_net159;
 wire clknet_1_0__leaf_net159;
 wire clknet_1_1__leaf_net159;
 wire clknet_0_net157;
 wire clknet_1_0__leaf_net157;
 wire clknet_1_1__leaf_net157;
 wire clknet_0_net658;
 wire clknet_1_0__leaf_net658;
 wire clknet_1_1__leaf_net658;
 wire clknet_0_net245;
 wire clknet_1_0__leaf_net245;
 wire clknet_1_1__leaf_net245;
 wire clknet_0_net657;
 wire clknet_1_0__leaf_net657;
 wire clknet_1_1__leaf_net657;
 wire clknet_0_net219;
 wire clknet_1_0__leaf_net219;
 wire clknet_1_1__leaf_net219;
 wire clknet_0_net231;
 wire clknet_1_0__leaf_net231;
 wire clknet_1_1__leaf_net231;
 wire clknet_0_net223;
 wire clknet_1_0__leaf_net223;
 wire clknet_1_1__leaf_net223;
 wire clknet_0_net229;
 wire clknet_1_0__leaf_net229;
 wire clknet_1_1__leaf_net229;
 wire clknet_0_net228;
 wire clknet_1_0__leaf_net228;
 wire clknet_1_1__leaf_net228;
 wire clknet_0_net220;
 wire clknet_1_0__leaf_net220;
 wire clknet_1_1__leaf_net220;
 wire clknet_0_net337;
 wire clknet_1_0__leaf_net337;
 wire clknet_1_1__leaf_net337;
 wire clknet_0_net212;
 wire clknet_1_0__leaf_net212;
 wire clknet_1_1__leaf_net212;
 wire net336;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;

 sky130_fd_sc_hd__a2111o_4 c100 (.A1(net812),
    .A2(net783),
    .B1(net805),
    .C1(net811),
    .D1(net806),
    .X(net854));
 sky130_fd_sc_hd__o2111ai_4 c101 (.A1(net789),
    .A2(net854),
    .B1(net785),
    .C1(net783),
    .D1(net806),
    .Y(net0));
 sky130_fd_sc_hd__a2111oi_2 c102 (.A1(net802),
    .A2(net854),
    .B1(net811),
    .C1(net812),
    .D1(net796),
    .Y(net1));
 sky130_fd_sc_hd__o2111a_1 c103 (.A1(net808),
    .A2(net1),
    .B1(net809),
    .C1(net811),
    .D1(net786),
    .X(net836));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net786),
    .A1(net791),
    .A2(net800),
    .A3(net813),
    .S0(net801),
    .S1(net769),
    .X(net837));
 sky130_fd_sc_hd__o2111ai_2 c105 (.A1(net809),
    .A2(net739),
    .B1(net808),
    .C1(net790),
    .D1(net837),
    .Y(net2));
 sky130_fd_sc_hd__mux4_1 c106 (.A0(net778),
    .A1(net811),
    .A2(net919),
    .A3(net837),
    .S0(net808),
    .S1(net810),
    .X(net867));
 sky130_fd_sc_hd__mux4_2 c107 (.A0(net2),
    .A1(net837),
    .A2(net867),
    .A3(net809),
    .S0(net811),
    .S1(net807),
    .X(net871));
 sky130_fd_sc_hd__o2111ai_4 c108 (.A1(net807),
    .A2(net787),
    .B1(net871),
    .C1(net811),
    .D1(net779),
    .Y(net3));
 sky130_fd_sc_hd__a2111oi_1 c109 (.A1(net3),
    .A2(net804),
    .B1(net802),
    .C1(net2),
    .D1(net721),
    .Y(net4));
 sky130_fd_sc_hd__nand3_2 c122 (.A(net783),
    .B(net804),
    .C(net810),
    .Y(net868));
 sky130_fd_sc_hd__nor2_2 c123 (.A(net813),
    .B(net868),
    .Y(net5));
 sky130_fd_sc_hd__nor3_2 c124 (.A(net752),
    .B(net782),
    .C(net5),
    .Y(net874));
 sky130_fd_sc_hd__o2111a_1 c125 (.A1(net801),
    .A2(net837),
    .B1(net796),
    .C1(net806),
    .D1(net790),
    .X(net851));
 sky130_fd_sc_hd__or3_4 c126 (.A(net5),
    .B(net913),
    .C(net748),
    .X(net877));
 sky130_fd_sc_hd__or4bb_2 c127 (.A(net877),
    .B(net806),
    .C_N(net5),
    .D_N(net913),
    .X(net879));
 sky130_fd_sc_hd__a2111o_2 c128 (.A1(net5),
    .A2(net879),
    .B1(net813),
    .C1(net877),
    .D1(net913),
    .X(net880));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net868),
    .A1(net919),
    .A2(net879),
    .A3(net877),
    .S0(net5),
    .S1(net880),
    .X(net878));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net769),
    .A1(net724),
    .A2(net878),
    .A3(net880),
    .S0(net913),
    .S1(net877),
    .X(net881));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net880),
    .A1(net878),
    .A2(net851),
    .A3(net881),
    .S0(net877),
    .S1(net5),
    .X(net876));
 sky130_fd_sc_hd__or2_4 c132 (.A(net724),
    .B(net770),
    .X(net6));
 sky130_fd_sc_hd__nor3b_4 c133 (.A(net761),
    .B(net720),
    .C_N(net927),
    .Y(net7));
 sky130_fd_sc_hd__nand2b_4 c134 (.A_N(net717),
    .B(net981),
    .Y(net8));
 sky130_fd_sc_hd__or4bb_4 c135 (.A(net751),
    .B(net981),
    .C_N(net927),
    .D_N(net8),
    .X(net9));
 sky130_fd_sc_hd__mux4_2 c136 (.A0(net720),
    .A1(net9),
    .A2(net8),
    .A3(net740),
    .S0(net981),
    .S1(net781),
    .X(net10));
 sky130_fd_sc_hd__or3_4 c137 (.A(net731),
    .B(net8),
    .C(net9),
    .X(net11));
 sky130_fd_sc_hd__or3b_4 c138 (.A(net792),
    .B(net7),
    .C_N(net909),
    .X(net12));
 sky130_fd_sc_hd__o2111ai_4 c139 (.A1(net727),
    .A2(net730),
    .B1(net770),
    .C1(net9),
    .D1(net725),
    .Y(net13));
 sky130_fd_sc_hd__o2111a_4 c140 (.A1(net981),
    .A2(net12),
    .B1(net929),
    .C1(net9),
    .D1(net719),
    .X(net14));
 sky130_fd_sc_hd__nand3b_4 c141 (.A_N(net8),
    .B(net14),
    .C(net717),
    .Y(net15));
 sky130_fd_sc_hd__and2b_2 c142 (.A_N(net781),
    .B(net717),
    .X(net16));
 sky130_fd_sc_hd__and2b_1 c143 (.A_N(net12),
    .B(net15),
    .X(net17));
 sky130_fd_sc_hd__or3b_4 c144 (.A(net16),
    .B(net726),
    .C_N(net17),
    .X(net18));
 sky130_fd_sc_hd__and3b_4 c145 (.A_N(net14),
    .B(net17),
    .C(net15),
    .X(net19));
 sky130_fd_sc_hd__nor3_4 c146 (.A(net724),
    .B(net16),
    .C(net18),
    .Y(net20));
 sky130_fd_sc_hd__o2111ai_4 c147 (.A1(net940),
    .A2(net740),
    .B1(net728),
    .C1(net15),
    .D1(net18),
    .Y(net21));
 sky130_fd_sc_hd__nor2b_1 c148 (.A(net21),
    .B_N(net717),
    .Y(net22));
 sky130_fd_sc_hd__a2111o_4 c149 (.A1(net20),
    .A2(net10),
    .B1(net981),
    .C1(net21),
    .D1(net12),
    .X(net23));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net17),
    .A1(net14),
    .A2(net22),
    .A3(net938),
    .S0(net986),
    .S1(net15),
    .X(net24));
 sky130_fd_sc_hd__or4bb_1 c151 (.A(net726),
    .B(net22),
    .C_N(net985),
    .D_N(net10),
    .X(net25));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net15),
    .A1(net986),
    .A2(net938),
    .A3(net22),
    .S0(net12),
    .S1(net909),
    .X(net873));
 sky130_fd_sc_hd__or4bb_1 c153 (.A(net990),
    .B(net986),
    .C_N(net22),
    .D_N(net873),
    .X(net26));
 sky130_fd_sc_hd__or2b_1 c154 (.A(net755),
    .B_N(net745),
    .X(net27));
 sky130_fd_sc_hd__or4bb_4 c155 (.A(net981),
    .B(net735),
    .C_N(net742),
    .D_N(net803),
    .X(net28));
 sky130_fd_sc_hd__nand2_1 c156 (.A(net14),
    .B(net770),
    .Y(net29));
 sky130_fd_sc_hd__nand3_1 c157 (.A(net733),
    .B(net747),
    .C(net918),
    .Y(net30));
 sky130_fd_sc_hd__or4bb_2 c158 (.A(net730),
    .B(net755),
    .C_N(net746),
    .D_N(net26),
    .X(net31));
 sky130_fd_sc_hd__and4b_4 c159 (.A_N(net746),
    .B(net29),
    .C(net739),
    .D(net9),
    .X(net32));
 sky130_fd_sc_hd__and2_4 c160 (.A(net745),
    .B(net30),
    .X(net33));
 sky130_fd_sc_hd__a2111o_2 c161 (.A1(net738),
    .A2(net13),
    .B1(net741),
    .C1(net770),
    .D1(net926),
    .X(net34));
 sky130_fd_sc_hd__nand2b_2 c162 (.A_N(net918),
    .B(net730),
    .Y(net35));
 sky130_fd_sc_hd__nor2_2 c163 (.A(net30),
    .B(net32),
    .Y(net36));
 sky130_fd_sc_hd__nand3_2 c164 (.A(net29),
    .B(net739),
    .C(net736),
    .Y(net37));
 sky130_fd_sc_hd__nor2_1 c165 (.A(net750),
    .B(net730),
    .Y(net872));
 sky130_fd_sc_hd__nor4b_1 c166 (.A(net741),
    .B(net755),
    .C(net754),
    .D_N(net918),
    .Y(net38));
 sky130_fd_sc_hd__nand3b_4 c167 (.A_N(net739),
    .B(net32),
    .C(net912),
    .Y(net39));
 sky130_fd_sc_hd__nor4b_2 c168 (.A(net39),
    .B(net9),
    .C(net749),
    .D_N(net735),
    .Y(net856));
 sky130_fd_sc_hd__or4_1 c169 (.A(net735),
    .B(net755),
    .C(net986),
    .D(net725),
    .X(net40));
 sky130_fd_sc_hd__a2111o_1 c170 (.A1(net40),
    .A2(net725),
    .B1(net872),
    .C1(net899),
    .D1(net926),
    .X(net41));
 sky130_fd_sc_hd__mux4_1 c171 (.A0(net27),
    .A1(net26),
    .A2(net30),
    .A3(net38),
    .S0(net32),
    .S1(net31),
    .X(net42));
 sky130_fd_sc_hd__or4b_1 c172 (.A(net42),
    .B(net36),
    .C(net747),
    .D_N(net746),
    .X(net43));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net34),
    .A1(net36),
    .A2(net42),
    .A3(net755),
    .S0(net742),
    .S1(net872),
    .X(net44));
 sky130_fd_sc_hd__a2111o_1 c174 (.A1(net856),
    .A2(net750),
    .B1(net41),
    .C1(net19),
    .D1(net626),
    .X(net45));
 sky130_fd_sc_hd__or4_1 c175 (.A(net33),
    .B(net42),
    .C(net32),
    .X(net46));
 sky130_fd_sc_hd__and3_1 c176 (.A(net766),
    .B(net747),
    .C(net734),
    .X(net47));
 sky130_fd_sc_hd__and3_2 c177 (.A(net26),
    .B(net39),
    .C(net626),
    .X(net864));
 sky130_fd_sc_hd__nor4b_2 c178 (.A(net775),
    .B(net24),
    .C(net35),
    .D_N(net626),
    .Y(net48));
 sky130_fd_sc_hd__a2111o_2 c179 (.A1(net754),
    .A2(net773),
    .B1(net927),
    .C1(net758),
    .D1(net924),
    .X(net49));
 sky130_fd_sc_hd__or4_1 c180 (.A(net736),
    .B(net758),
    .C(net33),
    .D(net756),
    .X(net50));
 sky130_fd_sc_hd__nor3b_2 c181 (.A(net768),
    .B(net49),
    .C_N(net924),
    .Y(net51));
 sky130_fd_sc_hd__nor3_1 c182 (.A(net756),
    .B(net759),
    .C(net924),
    .Y(net52));
 sky130_fd_sc_hd__nand3b_1 c183 (.A_N(net734),
    .B(net48),
    .C(net864),
    .Y(net53));
 sky130_fd_sc_hd__or3b_4 c184 (.A(net759),
    .B(net50),
    .C_N(net747),
    .X(net54));
 sky130_fd_sc_hd__nor3b_2 c185 (.A(net737),
    .B(net742),
    .C_N(net864),
    .Y(net55));
 sky130_fd_sc_hd__buf_6 c186 (.A(net620),
    .X(net56));
 sky130_fd_sc_hd__nand3_4 c187 (.A(net757),
    .B(net899),
    .C(net864),
    .Y(net859));
 sky130_fd_sc_hd__and4bb_1 c188 (.A_N(net864),
    .B_N(net52),
    .C(net763),
    .D(net35),
    .X(net57));
 sky130_fd_sc_hd__and4_1 c189 (.A(net911),
    .B(net54),
    .C(net24),
    .D(net864),
    .X(net58));
 sky130_fd_sc_hd__nor4_1 c190 (.A(net859),
    .B(net57),
    .C(net56),
    .D(net49),
    .Y(net59));
 sky130_fd_sc_hd__inv_1 c191 (.A(net620),
    .Y(net60));
 sky130_fd_sc_hd__inv_2 c192 (.A(net603),
    .Y(net61));
 sky130_fd_sc_hd__mux4_1 c193 (.A0(net772),
    .A1(net864),
    .A2(net58),
    .A3(net859),
    .S0(net773),
    .S1(net760),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net774),
    .A1(net54),
    .A2(net56),
    .A3(net60),
    .S0(net924),
    .S1(net603),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net764),
    .A1(net759),
    .A2(net48),
    .A3(net54),
    .S0(net872),
    .S1(net924),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 c196 (.A(net603),
    .X(net65));
 sky130_fd_sc_hd__mux4_2 c197 (.A0(net50),
    .A1(net64),
    .A2(net49),
    .A3(net65),
    .S0(net911),
    .S1(net754),
    .X(net66));
 sky130_fd_sc_hd__or3_2 c198 (.A(net788),
    .B(net924),
    .C(net603),
    .X(net67));
 sky130_fd_sc_hd__nand3b_4 c199 (.A_N(net60),
    .B(net788),
    .C(net67),
    .Y(net849));
 sky130_fd_sc_hd__or3_4 c200 (.A(net849),
    .B(net797),
    .C(net795),
    .X(net68));
 sky130_fd_sc_hd__nand3b_1 c201 (.A_N(net777),
    .B(net68),
    .C(net19),
    .Y(net69));
 sky130_fd_sc_hd__nor3b_2 c202 (.A(net797),
    .B(net36),
    .C_N(net68),
    .Y(net70));
 sky130_fd_sc_hd__nand3b_1 c203 (.A_N(net987),
    .B(net68),
    .C(net978),
    .Y(net71));
 sky130_fd_sc_hd__and3_1 c204 (.A(net68),
    .B(net49),
    .C(net780),
    .X(net72));
 sky130_fd_sc_hd__mux4_2 c205 (.A0(net49),
    .A1(net68),
    .A2(net60),
    .A3(net72),
    .S0(net917),
    .S1(net986),
    .X(net862));
 sky130_fd_sc_hd__nand3b_2 c206 (.A_N(net69),
    .B(net777),
    .C(net72),
    .Y(net863));
 sky130_fd_sc_hd__inv_4 c207 (.A(net609),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 c208 (.A(net609),
    .Y(net74));
 sky130_fd_sc_hd__and4bb_1 c209 (.A_N(net336),
    .B_N(net67),
    .C(net70),
    .D(net849),
    .X(net75));
 sky130_fd_sc_hd__or3_1 c210 (.A(net73),
    .B(net924),
    .C(net69),
    .X(net76));
 sky130_fd_sc_hd__mux4_1 c211 (.A0(net76),
    .A1(net849),
    .A2(net929),
    .A3(net935),
    .S0(net873),
    .S1(net55),
    .X(net77));
 sky130_fd_sc_hd__nor3b_2 c212 (.A(net71),
    .B(net798),
    .C_N(net76),
    .Y(net78));
 sky130_fd_sc_hd__or4_1 c213 (.A(net75),
    .B(net800),
    .C(net71),
    .D(net933),
    .X(net79));
 sky130_fd_sc_hd__mux4_4 c214 (.A0(net79),
    .A1(net929),
    .A2(net725),
    .A3(net799),
    .S0(net73),
    .S1(net652),
    .X(net80));
 sky130_fd_sc_hd__mux4_2 c215 (.A0(net74),
    .A1(net863),
    .A2(net36),
    .A3(net76),
    .S0(net862),
    .S1(net608),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net79),
    .A1(net68),
    .A2(net81),
    .A3(net74),
    .S0(net78),
    .S1(net609),
    .X(net82));
 sky130_fd_sc_hd__and4_1 c217 (.A(net67),
    .B(net81),
    .C(net721),
    .D(net863),
    .X(net83));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net771),
    .A1(net68),
    .A2(net79),
    .A3(net770),
    .S0(net75),
    .S1(net83),
    .X(net84));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net72),
    .A1(net67),
    .A2(net79),
    .A3(net336),
    .S0(net608),
    .S1(net652),
    .X(net85));
 sky130_fd_sc_hd__or2b_1 c220 (.A(net980),
    .B_N(net739),
    .X(net86));
 sky130_fd_sc_hd__nand2_1 c221 (.A(net805),
    .B(net621),
    .Y(net87));
 sky130_fd_sc_hd__or2b_1 c222 (.A(net87),
    .B_N(net86),
    .X(net88));
 sky130_fd_sc_hd__or4_1 c223 (.A(net86),
    .B(net859),
    .C(net904),
    .D(net621),
    .X(net89));
 sky130_fd_sc_hd__or2_1 c224 (.A(net86),
    .B(net621),
    .X(net90));
 sky130_fd_sc_hd__or2_4 c225 (.A(net805),
    .B(net871),
    .X(net91));
 sky130_fd_sc_hd__or2_4 c226 (.A(net90),
    .B(net88),
    .X(net829));
 sky130_fd_sc_hd__o2111a_4 c227 (.A1(net917),
    .A2(net811),
    .B1(net909),
    .C1(net794),
    .D1(net620),
    .X(net92));
 sky130_fd_sc_hd__and2_1 c228 (.A(net744),
    .B(net626),
    .X(net93));
 sky130_fd_sc_hd__a2111oi_4 c229 (.A1(net92),
    .A2(net91),
    .B1(net88),
    .C1(net904),
    .D1(net68),
    .Y(net860));
 sky130_fd_sc_hd__and2b_1 c230 (.A_N(net83),
    .B(net91),
    .X(net94));
 sky130_fd_sc_hd__nor2b_1 c231 (.A(net901),
    .B_N(net854),
    .Y(net95));
 sky130_fd_sc_hd__or3_4 c232 (.A(net95),
    .B(net873),
    .C(net93),
    .X(net96));
 sky130_fd_sc_hd__buf_6 c233 (.A(net621),
    .X(net97));
 sky130_fd_sc_hd__a2111oi_1 c234 (.A1(net94),
    .A2(net91),
    .B1(net3),
    .C1(net96),
    .D1(net860),
    .Y(net98));
 sky130_fd_sc_hd__a2111o_2 c235 (.A1(net836),
    .A2(net782),
    .B1(net90),
    .C1(net620),
    .D1(net621),
    .X(net861));
 sky130_fd_sc_hd__or2_4 c236 (.A(net861),
    .B(net621),
    .X(net99));
 sky130_fd_sc_hd__nor3b_1 c237 (.A(net93),
    .B(net87),
    .C_N(net901),
    .Y(net100));
 sky130_fd_sc_hd__or4_4 c238 (.A(net100),
    .B(net96),
    .C(net99),
    .D(net83),
    .X(net866));
 sky130_fd_sc_hd__mux4_2 c239 (.A0(net99),
    .A1(net100),
    .A2(net95),
    .A3(net3),
    .S0(net97),
    .S1(net849),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net36),
    .A1(net94),
    .A2(net866),
    .A3(net100),
    .S0(net96),
    .S1(net91),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net101),
    .A1(net100),
    .A2(net784),
    .A3(net99),
    .S0(net620),
    .S1(net621),
    .X(net870));
 sky130_fd_sc_hd__nand2b_2 c264 (.A_N(net723),
    .B(net19),
    .Y(net103));
 sky130_fd_sc_hd__nand3_4 c265 (.A(net740),
    .B(net929),
    .C(net770),
    .Y(net104));
 sky130_fd_sc_hd__and3b_2 c266 (.A_N(net719),
    .B(net19),
    .C(net929),
    .X(net105));
 sky130_fd_sc_hd__nand3_2 c267 (.A(net984),
    .B(net16),
    .C(net104),
    .Y(net106));
 sky130_fd_sc_hd__or3_1 c268 (.A(net25),
    .B(net103),
    .C(net22),
    .X(net107));
 sky130_fd_sc_hd__nor3_2 c269 (.A(net8),
    .B(net104),
    .C(net895),
    .Y(net108));
 sky130_fd_sc_hd__or3b_4 c270 (.A(net105),
    .B(net12),
    .C_N(net895),
    .X(net109));
 sky130_fd_sc_hd__or4_1 c271 (.A(net909),
    .B(net719),
    .C(net108),
    .D(net106),
    .X(net110));
 sky130_fd_sc_hd__or4b_1 c272 (.A(net22),
    .B(net21),
    .C(net15),
    .D_N(net885),
    .X(net111));
 sky130_fd_sc_hd__sdfbbn_2 c273 (.CLK_N(clknet_4_1_0_clk),
    .D(net15),
    .RESET_B(net12),
    .SCD(net895),
    .SCE(net885),
    .SET_B(net585),
    .Q(net113),
    .Q_N(net112));
 sky130_fd_sc_hd__sdfrbp_2 c274 (.CLK(clknet_4_4_0_clk),
    .D(net108),
    .RESET_B(net112),
    .SCD(net885),
    .SCE(net585),
    .Q(net115),
    .Q_N(net114));
 sky130_fd_sc_hd__dfbbn_1 c275 (.CLK_N(clknet_4_0_0_clk),
    .D(net115),
    .RESET_B(net723),
    .SET_B(net885),
    .Q(net117),
    .Q_N(net116));
 sky130_fd_sc_hd__sdfrbp_2 c276 (.CLK(clknet_4_1_0_clk),
    .D(net117),
    .RESET_B(net103),
    .SCD(net885),
    .SCE(net585),
    .Q(net119),
    .Q_N(net118));
 sky130_fd_sc_hd__nand3b_4 c277 (.A_N(net119),
    .B(net895),
    .C(net114),
    .Y(net852));
 sky130_fd_sc_hd__mux4_1 c278 (.A0(net103),
    .A1(net116),
    .A2(net885),
    .A3(net104),
    .S0(net852),
    .S1(net895),
    .X(net120));
 sky130_fd_sc_hd__or3b_2 c279 (.A(net895),
    .B(net103),
    .C_N(net104),
    .X(net121));
 sky130_fd_sc_hd__mux4_1 c280 (.A0(net852),
    .A1(net16),
    .A2(net121),
    .A3(net885),
    .S0(net895),
    .S1(net114),
    .X(net122));
 sky130_fd_sc_hd__sdfbbn_1 c281 (.CLK_N(clknet_4_1_0_clk),
    .D(net121),
    .RESET_B(net852),
    .SCD(net103),
    .SCE(net885),
    .SET_B(net655),
    .Q(net124),
    .Q_N(net123));
 sky130_fd_sc_hd__mux4_2 c282 (.A0(net121),
    .A1(net106),
    .A2(net124),
    .A3(net108),
    .S0(net852),
    .S1(net655),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net125),
    .A1(net124),
    .A2(net115),
    .A3(net108),
    .S0(net104),
    .S1(net585),
    .X(net126));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net121),
    .A1(net16),
    .A2(net123),
    .A3(net104),
    .S0(net885),
    .S1(net585),
    .X(net127));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net953),
    .A1(net121),
    .A2(net109),
    .A3(net125),
    .S0(net855),
    .S1(net656),
    .X(net128));
 sky130_fd_sc_hd__nor3_1 c286 (.A(net45),
    .B(net749),
    .C(net109),
    .Y(net129));
 sky130_fd_sc_hd__nand3b_2 c287 (.A_N(net912),
    .B(net938),
    .C(net749),
    .Y(net130));
 sky130_fd_sc_hd__nor3b_2 c288 (.A(net115),
    .B(net626),
    .C_N(net656),
    .Y(net131));
 sky130_fd_sc_hd__and3b_4 c289 (.A_N(net803),
    .B(net24),
    .C(net732),
    .X(net132));
 sky130_fd_sc_hd__nor3b_1 c290 (.A(net37),
    .B(net912),
    .C_N(net132),
    .Y(net133));
 sky130_fd_sc_hd__clkbuf_2 c291 (.A(net606),
    .X(net134));
 sky130_fd_sc_hd__and3b_1 c292 (.A_N(net131),
    .B(net45),
    .C(net626),
    .X(net135));
 sky130_fd_sc_hd__nand3b_2 c293 (.A_N(net32),
    .B(net134),
    .C(net131),
    .Y(net136));
 sky130_fd_sc_hd__mux4_2 c294 (.A0(net108),
    .A1(net724),
    .A2(net856),
    .A3(net132),
    .S0(net31),
    .S1(net655),
    .X(net137));
 sky130_fd_sc_hd__a2111oi_1 c295 (.A1(net31),
    .A2(net952),
    .B1(net131),
    .C1(net114),
    .D1(net112),
    .Y(net138));
 sky130_fd_sc_hd__inv_4 c296 (.A(net606),
    .Y(net139));
 sky130_fd_sc_hd__and4_1 c297 (.A(net136),
    .B(net133),
    .C(net139),
    .D(net134),
    .X(net140));
 sky130_fd_sc_hd__nand3b_2 c298 (.A_N(net103),
    .B(net32),
    .C(net656),
    .Y(net141));
 sky130_fd_sc_hd__nand3b_4 c299 (.A_N(net132),
    .B(net141),
    .C(net753),
    .Y(net142));
 sky130_fd_sc_hd__mux4_4 c300 (.A0(net133),
    .A1(net19),
    .A2(net743),
    .A3(net753),
    .S0(net886),
    .S1(net892),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 c301 (.A0(net13),
    .A1(net141),
    .A2(net134),
    .A3(net108),
    .S0(net129),
    .S1(net135),
    .X(net144));
 sky130_fd_sc_hd__sdfbbp_1 c302 (.CLK(clknet_4_4_0_clk),
    .D(net139),
    .RESET_B(net13),
    .SCD(net140),
    .SCE(net892),
    .SET_B(clknet_1_1__leaf_net658),
    .Q(net146),
    .Q_N(net145));
 sky130_fd_sc_hd__mux4_4 c303 (.A0(net131),
    .A1(net129),
    .A2(net977),
    .A3(net13),
    .S0(net132),
    .S1(clknet_1_0__leaf_net658),
    .X(net147));
 sky130_fd_sc_hd__mux4_2 c304 (.A0(net135),
    .A1(net136),
    .A2(net133),
    .A3(net137),
    .S0(net892),
    .S1(clknet_1_0__leaf_net658),
    .X(net148));
 sky130_fd_sc_hd__mux4_2 c305 (.A0(net140),
    .A1(net918),
    .A2(net130),
    .A3(clknet_1_1__leaf_net625),
    .S0(clknet_1_0__leaf_net658),
    .S1(clknet_1_0__leaf_net659),
    .X(net149));
 sky130_fd_sc_hd__mux4_2 c306 (.A0(net41),
    .A1(net134),
    .A2(net747),
    .A3(net605),
    .S0(clknet_1_0__leaf_net625),
    .S1(clknet_1_0__leaf_net659),
    .X(net150));
 sky130_fd_sc_hd__a2111o_2 c307 (.A1(clknet_1_0__leaf_net150),
    .A2(net139),
    .B1(net145),
    .C1(net605),
    .D1(clknet_1_0__leaf_net625),
    .X(net151));
 sky130_fd_sc_hd__or3b_1 c308 (.A(net63),
    .B(net35),
    .C_N(net893),
    .X(net152));
 sky130_fd_sc_hd__nand3_4 c309 (.A(net61),
    .B(net758),
    .C(net911),
    .Y(net153));
 sky130_fd_sc_hd__or4_2 c310 (.A(net747),
    .B(net119),
    .C(net24),
    .D(clknet_1_0__leaf_net659),
    .X(net154));
 sky130_fd_sc_hd__or3_2 c311 (.A(net776),
    .B(net65),
    .C(net928),
    .X(net155));
 sky130_fd_sc_hd__or3b_4 c312 (.A(clknet_1_1__leaf_net150),
    .B(net852),
    .C_N(net753),
    .X(net156));
 sky130_fd_sc_hd__nor3_1 c313 (.A(net65),
    .B(net908),
    .C(clknet_1_1__leaf_net154),
    .Y(net157));
 sky130_fd_sc_hd__inv_4 c314 (.A(net622),
    .Y(net158));
 sky130_fd_sc_hd__nand4_1 c315 (.A(net770),
    .B(clknet_1_0__leaf_net154),
    .C(net892),
    .D(net656),
    .Y(net159));
 sky130_fd_sc_hd__mux4_4 c316 (.A0(net106),
    .A1(net113),
    .A2(net152),
    .A3(clknet_1_0__leaf_net157),
    .S0(net893),
    .S1(clknet_1_0__leaf_net154),
    .X(net160));
 sky130_fd_sc_hd__nand3_2 c317 (.A(net35),
    .B(net132),
    .C(clknet_1_0__leaf_net154),
    .Y(net161));
 sky130_fd_sc_hd__nand4_1 c318 (.A(net897),
    .B(net145),
    .C(net892),
    .D(net638),
    .Y(net162));
 sky130_fd_sc_hd__inv_4 c319 (.A(net622),
    .Y(net163));
 sky130_fd_sc_hd__and4_2 c320 (.A(net163),
    .B(net158),
    .C(net908),
    .D(net893),
    .X(net164));
 sky130_fd_sc_hd__inv_1 c321 (.A(net623),
    .Y(net831));
 sky130_fd_sc_hd__or3_2 c322 (.A(net158),
    .B(clknet_1_0__leaf_net154),
    .C(clknet_1_0__leaf_net659),
    .X(net165));
 sky130_fd_sc_hd__sdfrtn_1 c323 (.CLK_N(clknet_4_5_0_clk),
    .D(net57),
    .RESET_B(net155),
    .SCD(net163),
    .SCE(net152),
    .Q(net166));
 sky130_fd_sc_hd__mux4_2 c324 (.A0(net753),
    .A1(clknet_1_0__leaf_net150),
    .A2(net923),
    .A3(clknet_1_0__leaf_net165),
    .S0(net145),
    .S1(net908),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net64),
    .A1(clknet_1_1__leaf_net150),
    .A2(net859),
    .A3(net33),
    .S0(net923),
    .S1(clknet_1_0__leaf_net659),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(clknet_1_0__leaf_net165),
    .A1(clknet_1_0__leaf_net159),
    .A2(net724),
    .A3(net158),
    .S0(net112),
    .S1(net923),
    .X(net169));
 sky130_fd_sc_hd__mux4_2 c327 (.A0(clknet_1_0__leaf_net167),
    .A1(net923),
    .A2(net724),
    .A3(net626),
    .S0(net644),
    .S1(net846),
    .X(net170));
 sky130_fd_sc_hd__mux4_2 c328 (.A0(clknet_1_0__leaf_net154),
    .A1(net61),
    .A2(net166),
    .A3(net908),
    .S0(net164),
    .S1(clknet_1_0__leaf_net625),
    .X(net171));
 sky130_fd_sc_hd__mux4_4 c329 (.A0(net166),
    .A1(net883),
    .A2(net65),
    .A3(net54),
    .S0(clknet_1_0__leaf_net161),
    .S1(net846),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 c330 (.A(net621),
    .X(net173));
 sky130_fd_sc_hd__nor3b_1 c331 (.A(net798),
    .B(net749),
    .C_N(net661),
    .Y(net174));
 sky130_fd_sc_hd__and4bb_1 c332 (.A_N(net78),
    .B_N(net142),
    .C(net626),
    .D(net964),
    .X(net175));
 sky130_fd_sc_hd__or3_4 c333 (.A(net70),
    .B(net173),
    .C(net661),
    .X(net176));
 sky130_fd_sc_hd__or3_2 c334 (.A(net174),
    .B(net893),
    .C(net626),
    .X(net177));
 sky130_fd_sc_hd__nor3b_2 c335 (.A(net780),
    .B(net779),
    .C_N(net846),
    .Y(net178));
 sky130_fd_sc_hd__nand3b_2 c336 (.A_N(net178),
    .B(net770),
    .C(net626),
    .Y(net179));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(net146),
    .A1(net19),
    .A2(net888),
    .A3(net70),
    .S0(net654),
    .S1(net855),
    .X(net180));
 sky130_fd_sc_hd__mux4_2 c338 (.A0(net176),
    .A1(net81),
    .A2(net760),
    .A3(net179),
    .S0(net603),
    .S1(net662),
    .X(net181));
 sky130_fd_sc_hd__a2111oi_0 c339 (.A1(net795),
    .A2(net908),
    .B1(net118),
    .C1(clknet_1_1__leaf_net659),
    .D1(net662),
    .Y(net182));
 sky130_fd_sc_hd__or4_4 c340 (.A(net916),
    .B(net791),
    .C(clknet_1_0__leaf_net182),
    .D(net663),
    .X(net183));
 sky130_fd_sc_hd__nor3b_2 c341 (.A(clknet_1_0__leaf_net182),
    .B(net916),
    .C_N(net660),
    .Y(net184));
 sky130_fd_sc_hd__mux4_2 c342 (.A0(net81),
    .A1(net780),
    .A2(net176),
    .A3(net652),
    .S0(net661),
    .S1(net662),
    .X(net838));
 sky130_fd_sc_hd__mux4_4 c343 (.A0(net799),
    .A1(net181),
    .A2(net70),
    .A3(clknet_1_0__leaf_net183),
    .S0(net164),
    .S1(clknet_1_0__leaf_net182),
    .X(net185));
 sky130_fd_sc_hd__mux4_4 c344 (.A0(clknet_1_1__leaf_net183),
    .A1(net178),
    .A2(net177),
    .A3(clknet_1_0__leaf_net182),
    .S0(net181),
    .S1(net660),
    .X(net186));
 sky130_fd_sc_hd__a2111o_2 c345 (.A1(net19),
    .A2(net178),
    .B1(net181),
    .C1(clknet_1_0__leaf_net182),
    .D1(net663),
    .X(net844));
 sky130_fd_sc_hd__mux4_2 c346 (.A0(net78),
    .A1(net181),
    .A2(net779),
    .A3(clknet_1_0__leaf_net844),
    .S0(net179),
    .S1(clknet_1_0__leaf_net182),
    .X(net187));
 sky130_fd_sc_hd__mux4_2 c347 (.A0(net173),
    .A1(net179),
    .A2(clknet_1_0__leaf_net183),
    .A3(clknet_1_0__leaf_net154),
    .S0(clknet_1_0__leaf_net844),
    .S1(net664),
    .X(net188));
 sky130_fd_sc_hd__and4_4 c348 (.A(net164),
    .B(clknet_1_0__leaf_net844),
    .C(clknet_1_0__leaf_net182),
    .D(net847),
    .X(net189));
 sky130_fd_sc_hd__a2111o_2 c349 (.A1(net70),
    .A2(net176),
    .B1(clknet_1_0__leaf_net182),
    .C1(clknet_1_0__leaf_net184),
    .D1(net888),
    .X(net190));
 sky130_fd_sc_hd__mux4_2 c350 (.A0(net849),
    .A1(net582),
    .A2(net638),
    .A3(net839),
    .S0(net663),
    .S1(net827),
    .X(net853));
 sky130_fd_sc_hd__mux4_4 c351 (.A0(clknet_1_0__leaf_net182),
    .A1(net853),
    .A2(net955),
    .A3(net582),
    .S0(net846),
    .S1(clknet_1_1__leaf_net659),
    .X(net191));
 sky130_fd_sc_hd__o2111ai_4 c352 (.A1(net804),
    .A2(net900),
    .B1(clknet_1_0__leaf_net182),
    .C1(net846),
    .D1(net827),
    .Y(net192));
 sky130_fd_sc_hd__a2111o_1 c353 (.A1(net97),
    .A2(net92),
    .B1(net794),
    .C1(net804),
    .D1(net893),
    .X(net193));
 sky130_fd_sc_hd__a2111oi_1 c354 (.A1(net760),
    .A2(net836),
    .B1(net926),
    .C1(net893),
    .D1(net855),
    .Y(net194));
 sky130_fd_sc_hd__a2111oi_4 c355 (.A1(net0),
    .A2(net132),
    .B1(net935),
    .C1(net782),
    .D1(clknet_1_0__leaf_net182),
    .Y(net195));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net882),
    .A1(net793),
    .A2(net861),
    .A3(net101),
    .S0(net99),
    .S1(net848),
    .X(net196));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net770),
    .A1(net811),
    .A2(net909),
    .A3(net782),
    .S0(net3),
    .S1(net610),
    .X(net197));
 sky130_fd_sc_hd__mux4_2 c358 (.A0(net193),
    .A1(net898),
    .A2(net0),
    .A3(net744),
    .S0(clknet_1_1__leaf_net192),
    .S1(net91),
    .X(net198));
 sky130_fd_sc_hd__mux4_2 c359 (.A0(clknet_1_1__leaf_net192),
    .A1(net97),
    .A2(clknet_1_0__leaf_net195),
    .A3(net936),
    .S0(net610),
    .S1(net847),
    .X(net199));
 sky130_fd_sc_hd__mux4_2 c360 (.A0(net199),
    .A1(net101),
    .A2(net3),
    .A3(net866),
    .S0(net193),
    .S1(net651),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net197),
    .A1(net785),
    .A2(net900),
    .A3(net853),
    .S0(net92),
    .S1(net804),
    .X(net845));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(net97),
    .A1(net51),
    .A2(net882),
    .A3(net924),
    .S0(net894),
    .S1(net651),
    .X(net201));
 sky130_fd_sc_hd__mux4_2 c363 (.A0(net849),
    .A1(net197),
    .A2(net101),
    .A3(net852),
    .S0(net581),
    .S1(net635),
    .X(net843));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net191),
    .A1(net838),
    .A2(net901),
    .A3(clknet_1_0__leaf_net192),
    .S0(net852),
    .S1(net652),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net794),
    .A1(clknet_1_0__leaf_net192),
    .A2(net859),
    .A3(net101),
    .S0(net742),
    .S1(net581),
    .X(net203));
 sky130_fd_sc_hd__nor4b_1 c366 (.A(net935),
    .B(net782),
    .C(clknet_1_0__leaf_net202),
    .D_N(net582),
    .Y(net204));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net132),
    .A1(clknet_1_0__leaf_net156),
    .A2(net852),
    .A3(net843),
    .S0(net847),
    .S1(net848),
    .X(net205));
 sky130_fd_sc_hd__a2111oi_2 c368 (.A1(net181),
    .A2(net51),
    .B1(net758),
    .C1(net724),
    .D1(clknet_1_0__leaf_net182),
    .Y(net206));
 sky130_fd_sc_hd__mux4_2 c369 (.A0(clknet_1_1__leaf_net157),
    .A1(net3),
    .A2(net843),
    .A3(net854),
    .S0(clknet_1_0__leaf_net206),
    .S1(net651),
    .X(net207));
 sky130_fd_sc_hd__mux4_2 c370 (.A0(clknet_1_1__leaf_net202),
    .A1(net861),
    .A2(net937),
    .A3(net651),
    .S0(net848),
    .S1(net666),
    .X(net208));
 sky130_fd_sc_hd__o2111a_2 c371 (.A1(clknet_1_1__leaf_net206),
    .A2(net132),
    .B1(net849),
    .C1(net842),
    .D1(net666),
    .X(net209));
 sky130_fd_sc_hd__mux4_4 c372 (.A0(net800),
    .A1(net0),
    .A2(net635),
    .A3(net847),
    .S0(net842),
    .S1(net666),
    .X(net857));
 sky130_fd_sc_hd__a2111o_1 c373 (.A1(net843),
    .A2(net724),
    .B1(net770),
    .C1(net847),
    .D1(net666),
    .X(net210));
 sky130_fd_sc_hd__and2_1 c396 (.A(net104),
    .B(net728),
    .X(net211));
 sky130_fd_sc_hd__or4b_2 c397 (.A(net109),
    .B(net117),
    .C(net105),
    .D_N(clknet_1_0__leaf_net657),
    .X(net212));
 sky130_fd_sc_hd__and2_1 c398 (.A(net211),
    .B(net107),
    .X(net213));
 sky130_fd_sc_hd__nand3_4 c399 (.A(net20),
    .B(net118),
    .C(net929),
    .Y(net214));
 sky130_fd_sc_hd__clkbuf_2 c400 (.A(net961),
    .X(net215));
 sky130_fd_sc_hd__sdfbbn_1 c401 (.CLK_N(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net212),
    .RESET_B(net215),
    .SCD(net941),
    .SCE(net214),
    .SET_B(clknet_1_0__leaf_net657),
    .Q(net217),
    .Q_N(net216));
 sky130_fd_sc_hd__or3_4 c402 (.A(net215),
    .B(net118),
    .C(net214),
    .X(net218));
 sky130_fd_sc_hd__or3_4 c403 (.A(net740),
    .B(net214),
    .C(clknet_1_1__leaf_net657),
    .X(net219));
 sky130_fd_sc_hd__or3_2 c404 (.A(net124),
    .B(clknet_1_0__leaf_net219),
    .C(net218),
    .X(net220));
 sky130_fd_sc_hd__nand3b_1 c405 (.A_N(net16),
    .B(net214),
    .C(net215),
    .Y(net221));
 sky130_fd_sc_hd__and4bb_4 c406 (.A_N(net213),
    .B_N(net217),
    .C(net105),
    .D(net214),
    .X(net222));
 sky130_fd_sc_hd__nand3b_2 c407 (.A_N(net221),
    .B(clknet_1_1__leaf_net219),
    .C(clknet_1_0__leaf_net220),
    .Y(net223));
 sky130_fd_sc_hd__sdfbbn_2 c408 (.CLK_N(clknet_4_0_0_clk),
    .D(net214),
    .RESET_B(clknet_1_1__leaf_net212),
    .SCD(net213),
    .SCE(clknet_1_0__leaf_net220),
    .SET_B(net215),
    .Q(net225),
    .Q_N(net224));
 sky130_fd_sc_hd__sdfbbp_1 c409 (.CLK(clknet_4_0_0_clk),
    .D(net104),
    .RESET_B(net215),
    .SCD(net216),
    .SCE(net222),
    .SET_B(net975),
    .Q(net227),
    .Q_N(net226));
 sky130_fd_sc_hd__and3b_1 c410 (.A_N(clknet_1_0__leaf_net223),
    .B(net225),
    .C(net226),
    .X(net228));
 sky130_fd_sc_hd__or3b_2 c411 (.A(net215),
    .B(net25),
    .C_N(clknet_1_1__leaf_net223),
    .X(net229));
 sky130_fd_sc_hd__sdfrtp_1 c412 (.CLK(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net229),
    .RESET_B(net211),
    .SCD(net226),
    .SCE(net123),
    .Q(net230));
 sky130_fd_sc_hd__nand3_1 c413 (.A(clknet_1_0__leaf_net219),
    .B(clknet_1_0__leaf_net223),
    .C(clknet_1_0__leaf_net220),
    .Y(net231));
 sky130_fd_sc_hd__mux4_4 c414 (.A0(net10),
    .A1(net230),
    .A2(net116),
    .A3(net215),
    .S0(net222),
    .S1(net728),
    .X(net232));
 sky130_fd_sc_hd__inv_2 c415 (.A(net961),
    .Y(net233));
 sky130_fd_sc_hd__mux4_2 c416 (.A0(net233),
    .A1(net222),
    .A2(net230),
    .A3(clknet_1_0__leaf_net212),
    .S0(net942),
    .S1(net667),
    .X(net234));
 sky130_fd_sc_hd__mux4_4 c417 (.A0(net230),
    .A1(net105),
    .A2(net233),
    .A3(clknet_1_1__leaf_net229),
    .S0(clknet_1_0__leaf_net228),
    .S1(net16),
    .X(net235));
 sky130_fd_sc_hd__or3b_2 c418 (.A(net134),
    .B(net37),
    .C_N(net892),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 c419 (.A(net616),
    .X(net237));
 sky130_fd_sc_hd__clkinv_4 c420 (.A(net632),
    .Y(net238));
 sky130_fd_sc_hd__or3b_4 c421 (.A(net237),
    .B(net39),
    .C_N(net130),
    .X(net239));
 sky130_fd_sc_hd__nor2b_1 c422 (.A(net239),
    .B_N(net237),
    .Y(net240));
 sky130_fd_sc_hd__or2_1 c423 (.A(net240),
    .B(net113),
    .X(net241));
 sky130_fd_sc_hd__nand2_2 c424 (.A(net241),
    .B(net606),
    .Y(net242));
 sky130_fd_sc_hd__and3_2 c425 (.A(net926),
    .B(net227),
    .C(net242),
    .X(net243));
 sky130_fd_sc_hd__mux4_2 c426 (.A0(net241),
    .A1(net242),
    .A2(net953),
    .A3(net240),
    .S0(net222),
    .S1(clknet_1_0__leaf_net151),
    .X(net244));
 sky130_fd_sc_hd__or3b_4 c427 (.A(net892),
    .B(clknet_1_1__leaf_net658),
    .C_N(net669),
    .X(net245));
 sky130_fd_sc_hd__buf_6 c428 (.A(net616),
    .X(net246));
 sky130_fd_sc_hd__sdfrtp_4 c429 (.CLK(clknet_4_4_0_clk),
    .D(net141),
    .RESET_B(net242),
    .SCD(clknet_1_0__leaf_net245),
    .SCE(net892),
    .Q(net247));
 sky130_fd_sc_hd__clkbuf_2 c430 (.A(net616),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 c431 (.A(net616),
    .X(net249));
 sky130_fd_sc_hd__sdfbbn_1 c432 (.CLK_N(clknet_4_3_0_clk),
    .D(net222),
    .RESET_B(net225),
    .SCD(net249),
    .SCE(net247),
    .SET_B(clknet_1_1__leaf_net658),
    .Q(net251),
    .Q_N(net250));
 sky130_fd_sc_hd__a2111oi_0 c433 (.A1(net241),
    .A2(net242),
    .B1(clknet_1_1__leaf_net220),
    .C1(clknet_1_0__leaf_net151),
    .D1(net669),
    .Y(net252));
 sky130_fd_sc_hd__and3_1 c434 (.A(net249),
    .B(net600),
    .C(net669),
    .X(net253));
 sky130_fd_sc_hd__o2111a_1 c435 (.A1(net246),
    .A2(net109),
    .B1(net240),
    .C1(net892),
    .D1(net243),
    .X(net254));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net105),
    .A1(net37),
    .A2(net242),
    .A3(net249),
    .S0(net600),
    .S1(net669),
    .X(net255));
 sky130_fd_sc_hd__sdfbbn_2 c437 (.CLK_N(clknet_4_3_0_clk),
    .D(net249),
    .RESET_B(net253),
    .SCD(net255),
    .SCE(net939),
    .SET_B(net227),
    .Q(net257),
    .Q_N(net256));
 sky130_fd_sc_hd__mux4_2 c438 (.A0(net257),
    .A1(clknet_1_0__leaf_net245),
    .A2(net247),
    .A3(net249),
    .S0(net585),
    .S1(net669),
    .X(net258));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net253),
    .A1(net222),
    .A2(net247),
    .A3(net256),
    .S0(net893),
    .S1(net970),
    .X(net259));
 sky130_fd_sc_hd__buf_16 c440 (.A(net594),
    .X(net260));
 sky130_fd_sc_hd__nor3b_2 c441 (.A(net155),
    .B(net118),
    .C_N(net893),
    .Y(net261));
 sky130_fd_sc_hd__buf_1 c442 (.A(net593),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 c443 (.A(net631),
    .X(net263));
 sky130_fd_sc_hd__buf_2 c444 (.A(net629),
    .X(net264));
 sky130_fd_sc_hd__o2111a_1 c445 (.A1(net39),
    .A2(net744),
    .B1(net224),
    .C1(net264),
    .D1(net620),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(net264),
    .A1(net222),
    .A2(net883),
    .A3(net744),
    .S0(net831),
    .S1(net248),
    .X(net266));
 sky130_fd_sc_hd__nor3_1 c447 (.A(net260),
    .B(net248),
    .C(net264),
    .Y(net267));
 sky130_fd_sc_hd__nor4_2 c448 (.A(net260),
    .B(net247),
    .C(net262),
    .D(net638),
    .Y(net268));
 sky130_fd_sc_hd__inv_8 c449 (.A(net632),
    .Y(net269));
 sky130_fd_sc_hd__sdfrtp_1 c450 (.CLK(clknet_4_12_0_clk),
    .D(net268),
    .RESET_B(net963),
    .SCD(clknet_1_0__leaf_net245),
    .SCE(net594),
    .Q(net270));
 sky130_fd_sc_hd__or3_1 c451 (.A(net262),
    .B(net54),
    .C(net119),
    .X(net271));
 sky130_fd_sc_hd__or3b_1 c452 (.A(net218),
    .B(net270),
    .C_N(net617),
    .X(net272));
 sky130_fd_sc_hd__sdfsbp_1 c453 (.CLK(clknet_4_13_0_clk),
    .D(net271),
    .SCD(net264),
    .SCE(net908),
    .SET_B(net887),
    .Q(net274),
    .Q_N(net273));
 sky130_fd_sc_hd__sdfsbp_1 c454 (.CLK(clknet_4_12_0_clk),
    .D(net222),
    .SCD(net974),
    .SCE(net262),
    .SET_B(clknet_1_1__leaf_net231),
    .Q(net276),
    .Q_N(net275));
 sky130_fd_sc_hd__buf_4 c455 (.A(net629),
    .X(net277));
 sky130_fd_sc_hd__nor3_1 c456 (.A(net267),
    .B(net155),
    .C(net277),
    .Y(net278));
 sky130_fd_sc_hd__inv_4 c457 (.A(net623),
    .Y(net279));
 sky130_fd_sc_hd__nor3_1 c458 (.A(net272),
    .B(net907),
    .C(net894),
    .Y(net280));
 sky130_fd_sc_hd__mux4_4 c459 (.A0(net280),
    .A1(net279),
    .A2(net268),
    .A3(net275),
    .S0(net925),
    .S1(clknet_1_1__leaf_net165),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net270),
    .A1(net247),
    .A2(net279),
    .A3(net272),
    .S0(net261),
    .S1(net277),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net279),
    .A1(net991),
    .A2(net66),
    .A3(net278),
    .S0(net270),
    .S1(net260),
    .X(net283));
 sky130_fd_sc_hd__sdfstp_1 c462 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net184),
    .SCD(net177),
    .SCE(net238),
    .SET_B(clknet_1_1__leaf_net245),
    .Q(net284));
 sky130_fd_sc_hd__mux4_4 c463 (.A0(clknet_1_1__leaf_net184),
    .A1(net924),
    .A2(net238),
    .A3(net949),
    .S0(net638),
    .S1(net644),
    .X(net285));
 sky130_fd_sc_hd__nor3_2 c464 (.A(clknet_1_0__leaf_net285),
    .B(net894),
    .C(net670),
    .Y(net286));
 sky130_fd_sc_hd__nand4b_4 c465 (.A_N(net248),
    .B(clknet_1_0__leaf_net285),
    .C(clknet_1_1__leaf_net182),
    .D(net653),
    .Y(net287));
 sky130_fd_sc_hd__nand4b_1 c466 (.A_N(net274),
    .B(clknet_1_1__leaf_net184),
    .C(net894),
    .D(net673),
    .Y(net288));
 sky130_fd_sc_hd__mux4_2 c467 (.A0(net951),
    .A1(net284),
    .A2(net238),
    .A3(clknet_1_0__leaf_net288),
    .S0(clknet_1_1__leaf_net182),
    .S1(net653),
    .X(net289));
 sky130_fd_sc_hd__o2111ai_1 c468 (.A1(clknet_1_1__leaf_net287),
    .A2(clknet_1_0__leaf_net286),
    .B1(net929),
    .C1(net638),
    .D1(net674),
    .Y(net290));
 sky130_fd_sc_hd__sdfbbp_1 c469 (.CLK(clknet_4_13_0_clk),
    .D(net261),
    .RESET_B(clknet_1_1__leaf_net154),
    .SCD(net274),
    .SCE(net950),
    .SET_B(net664),
    .Q(net292),
    .Q_N(net291));
 sky130_fd_sc_hd__mux4_4 c470 (.A0(net276),
    .A1(net784),
    .A2(net888),
    .A3(net145),
    .S0(clknet_1_1__leaf_net286),
    .S1(net273),
    .X(net293));
 sky130_fd_sc_hd__o2111ai_2 c471 (.A1(clknet_1_0__leaf_net287),
    .A2(net800),
    .B1(net957),
    .C1(net749),
    .D1(clknet_1_1__leaf_net154),
    .Y(net294));
 sky130_fd_sc_hd__mux4_4 c472 (.A0(net178),
    .A1(clknet_1_0__leaf_net294),
    .A2(net887),
    .A3(net765),
    .S0(net673),
    .S1(net675),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net831),
    .A1(clknet_1_0__leaf_net184),
    .A2(net275),
    .A3(net33),
    .S0(net291),
    .S1(clknet_1_0__leaf_net676),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net292),
    .A1(net274),
    .A2(net749),
    .A3(clknet_1_1__leaf_net286),
    .S0(net277),
    .S1(net591),
    .X(net297));
 sky130_fd_sc_hd__mux4_4 c475 (.A0(clknet_1_1__leaf_net296),
    .A1(net276),
    .A2(net897),
    .A3(net894),
    .S0(net743),
    .S1(net273),
    .X(net298));
 sky130_fd_sc_hd__mux4_2 c476 (.A0(net284),
    .A1(net178),
    .A2(net910),
    .A3(clknet_1_1__leaf_net844),
    .S0(net675),
    .S1(clknet_1_1__leaf_net677),
    .X(net299));
 sky130_fd_sc_hd__mux4_4 c477 (.A0(clknet_1_1__leaf_net288),
    .A1(clknet_1_0__leaf_net296),
    .A2(net929),
    .A3(clknet_1_0__leaf_net294),
    .S0(clknet_1_0__leaf_net676),
    .S1(clknet_1_0__leaf_net678),
    .X(net300));
 sky130_fd_sc_hd__sdfbbn_2 c478 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net844),
    .RESET_B(net779),
    .SCD(net591),
    .SCE(clknet_1_1__leaf_net676),
    .SET_B(clknet_1_1__leaf_net677),
    .Q(net826),
    .Q_N(net301));
 sky130_fd_sc_hd__mux4_2 c479 (.A0(net119),
    .A1(net826),
    .A2(net249),
    .A3(net928),
    .S0(net922),
    .S1(clknet_1_1__leaf_net676),
    .X(net302));
 sky130_fd_sc_hd__sdfbbn_1 c480 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net286),
    .RESET_B(net301),
    .SCD(net675),
    .SCE(clknet_1_1__leaf_net676),
    .SET_B(clknet_1_1__leaf_net678),
    .Q(net304),
    .Q_N(net303));
 sky130_fd_sc_hd__a2111oi_1 c481 (.A1(net304),
    .A2(net910),
    .B1(net142),
    .C1(net591),
    .D1(clknet_1_0__leaf_net678),
    .Y(net305));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net302),
    .A1(net779),
    .A2(clknet_1_1__leaf_net305),
    .A3(net248),
    .S0(net301),
    .S1(clknet_1_1__leaf_net677),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net304),
    .A1(net153),
    .A2(net826),
    .A3(net291),
    .S0(clknet_1_0__leaf_net296),
    .S1(clknet_1_0__leaf_net302),
    .X(net307));
 sky130_fd_sc_hd__o2111a_2 c484 (.A1(net758),
    .A2(net811),
    .B1(net277),
    .C1(net894),
    .D1(net837),
    .X(net841));
 sky130_fd_sc_hd__sdfbbp_1 c485 (.CLK(clknet_4_15_0_clk),
    .D(net829),
    .RESET_B(net926),
    .SCD(net92),
    .SCE(net841),
    .SET_B(net680),
    .Q(net309),
    .Q_N(net308));
 sky130_fd_sc_hd__o2111ai_4 c486 (.A1(net888),
    .A2(net829),
    .B1(clknet_1_1__leaf_net285),
    .C1(clknet_1_1__leaf_net298),
    .D1(net91),
    .Y(net310));
 sky130_fd_sc_hd__mux4_2 c487 (.A0(net101),
    .A1(net91),
    .A2(clknet_1_0__leaf_net294),
    .A3(net92),
    .S0(clknet_1_1__leaf_net231),
    .S1(net834),
    .X(net311));
 sky130_fd_sc_hd__sdfbbn_2 c488 (.CLK_N(clknet_4_13_0_clk),
    .D(net309),
    .RESET_B(net866),
    .SCD(net758),
    .SCE(net34),
    .SET_B(net968),
    .Q(net313),
    .Q_N(net312));
 sky130_fd_sc_hd__mux4_2 c489 (.A0(net292),
    .A1(net99),
    .A2(net837),
    .A3(clknet_1_1__leaf_net182),
    .S0(net665),
    .S1(net828),
    .X(net314));
 sky130_fd_sc_hd__mux4_2 c490 (.A0(clknet_1_0__leaf_net307),
    .A1(net843),
    .A2(net990),
    .A3(clknet_1_0__leaf_net156),
    .S0(net929),
    .S1(net666),
    .X(net315));
 sky130_fd_sc_hd__mux4_2 c491 (.A0(clknet_1_0__leaf_net195),
    .A1(net838),
    .A2(net765),
    .A3(net101),
    .S0(net99),
    .S1(net665),
    .X(net316));
 sky130_fd_sc_hd__mux4_4 c492 (.A0(clknet_1_0__leaf_net314),
    .A1(net308),
    .A2(net811),
    .A3(net894),
    .S0(net830),
    .S1(net842),
    .X(net317));
 sky130_fd_sc_hd__mux4_2 c493 (.A0(net758),
    .A1(net837),
    .A2(clknet_1_1__leaf_net317),
    .A3(clknet_1_0__leaf_net307),
    .S0(net784),
    .S1(net635),
    .X(net318));
 sky130_fd_sc_hd__mux4_2 c494 (.A0(net959),
    .A1(clknet_1_1__leaf_net316),
    .A2(clknet_1_1__leaf_net314),
    .A3(net635),
    .S0(net665),
    .S1(net683),
    .X(net319));
 sky130_fd_sc_hd__mux4_4 c495 (.A0(clknet_1_1__leaf_net317),
    .A1(net313),
    .A2(net277),
    .A3(net837),
    .S0(net894),
    .S1(net666),
    .X(net320));
 sky130_fd_sc_hd__mux4_4 c496 (.A0(clknet_1_0__leaf_net317),
    .A1(net743),
    .A2(net92),
    .A3(clknet_1_1__leaf_net307),
    .S0(net681),
    .S1(net682),
    .X(net321));
 sky130_fd_sc_hd__mux4_2 c497 (.A0(clknet_1_0__leaf_net317),
    .A1(net309),
    .A2(net894),
    .A3(net673),
    .S0(net680),
    .S1(net684),
    .X(net322));
 sky130_fd_sc_hd__mux4_4 c498 (.A0(net101),
    .A1(clknet_1_1__leaf_net316),
    .A2(net785),
    .A3(net840),
    .S0(net683),
    .S1(net835),
    .X(net323));
 sky130_fd_sc_hd__mux4_2 c499 (.A0(clknet_1_1__leaf_net316),
    .A1(clknet_1_1__leaf_net195),
    .A2(net926),
    .A3(net665),
    .S0(net682),
    .S1(net684),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net894),
    .A1(clknet_1_1__leaf_net317),
    .A2(net679),
    .A3(net681),
    .S0(net850),
    .S1(net686),
    .X(net325));
 sky130_fd_sc_hd__mux4_2 c501 (.A0(clknet_1_1__leaf_net844),
    .A1(net829),
    .A2(clknet_1_1__leaf_net316),
    .A3(net784),
    .S0(net830),
    .S1(net686),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(clknet_1_1__leaf_net156),
    .A1(net833),
    .A2(net839),
    .A3(net684),
    .S0(net685),
    .S1(net686),
    .X(net327));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(clknet_1_1__leaf_net285),
    .A1(clknet_1_0__leaf_net317),
    .A2(net834),
    .A3(net684),
    .S0(net850),
    .S1(net686),
    .X(net328));
 sky130_fd_sc_hd__mux4_4 c504 (.A0(net779),
    .A1(net92),
    .A2(net308),
    .A3(net841),
    .S0(net834),
    .S1(net830),
    .X(net329));
 sky130_fd_sc_hd__mux4_2 c505 (.A0(net96),
    .A1(net820),
    .A2(net666),
    .A3(net684),
    .S0(net685),
    .S1(net686),
    .X(net819));
 sky130_fd_sc_hd__and3b_1 c528 (.A_N(net215),
    .B(net227),
    .C(net929),
    .X(net330));
 sky130_fd_sc_hd__nor3b_2 c529 (.A(net230),
    .B(net226),
    .C_N(net667),
    .Y(net331));
 sky130_fd_sc_hd__and3_1 c530 (.A(net330),
    .B(net109),
    .C(net915),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd1_1 c531 (.A(clknet_1_0__leaf_net714),
    .X(net333));
 sky130_fd_sc_hd__or2_2 c532 (.A(net915),
    .B(net728),
    .X(net334));
 sky130_fd_sc_hd__nand3_1 c533 (.A(net334),
    .B(net895),
    .C(net915),
    .Y(net335));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__o2111a_2 c535 (.A1(net221),
    .A2(net334),
    .B1(clknet_1_0__leaf_net220),
    .C1(net889),
    .D1(net667),
    .X(net337));
 sky130_fd_sc_hd__or4b_2 c536 (.A(clknet_1_1__leaf_net337),
    .B(clknet_1_0__leaf_net333),
    .C(net112),
    .D_N(net889),
    .X(net338));
 sky130_fd_sc_hd__clkinv_4 c537 (.A(net649),
    .Y(net339));
 sky130_fd_sc_hd__nand4b_4 c538 (.A_N(net728),
    .B(net339),
    .C(net334),
    .D(net889),
    .Y(net340));
 sky130_fd_sc_hd__nor4_1 c539 (.A(net895),
    .B(net340),
    .C(net891),
    .Y(net341));
 sky130_fd_sc_hd__or4b_1 c540 (.A(net213),
    .B(net339),
    .C(net227),
    .D_N(net889),
    .X(net342));
 sky130_fd_sc_hd__inv_6 c541 (.A(net649),
    .Y(net343));
 sky130_fd_sc_hd__mux4_1 c542 (.A0(net340),
    .A1(net218),
    .A2(net339),
    .A3(net334),
    .S0(net342),
    .S1(net343),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net339),
    .A1(net343),
    .A2(net340),
    .A3(clknet_1_1__leaf_net220),
    .S0(net334),
    .S1(net889),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net342),
    .A1(net340),
    .A2(net339),
    .A3(net343),
    .S0(net588),
    .S1(net689),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net340),
    .A1(net109),
    .A2(net339),
    .A3(net915),
    .S0(net588),
    .S1(net971),
    .X(net347));
 sky130_fd_sc_hd__mux4_4 c546 (.A0(net218),
    .A1(net340),
    .A2(net588),
    .A3(net615),
    .S0(net688),
    .S1(net690),
    .X(net348));
 sky130_fd_sc_hd__sdfbbn_1 c547 (.CLK_N(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net229),
    .RESET_B(net343),
    .SCD(net889),
    .SCE(net615),
    .SET_B(net690),
    .Q(net350),
    .Q_N(net349));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net332),
    .A1(net343),
    .A2(net895),
    .A3(net221),
    .S0(net339),
    .S1(net689),
    .X(net351));
 sky130_fd_sc_hd__a2111o_1 c549 (.A1(net117),
    .A2(net343),
    .B1(net889),
    .C1(net634),
    .D1(net648),
    .X(net352));
 sky130_fd_sc_hd__inv_6 c550 (.A(net580),
    .Y(net353));
 sky130_fd_sc_hd__inv_1 c551 (.A(net580),
    .Y(net354));
 sky130_fd_sc_hd__nor3b_4 c552 (.A(net246),
    .B(clknet_1_1__leaf_net333),
    .C_N(net918),
    .Y(net355));
 sky130_fd_sc_hd__sdfstp_2 c553 (.CLK(clknet_4_3_0_clk),
    .D(net125),
    .SCD(net928),
    .SCE(net249),
    .SET_B(net967),
    .Q(net356));
 sky130_fd_sc_hd__clkbuf_2 c554 (.A(net579),
    .X(net357));
 sky130_fd_sc_hd__and3_4 c555 (.A(net938),
    .B(net354),
    .C(net617),
    .X(net358));
 sky130_fd_sc_hd__nand4b_4 c556 (.A_N(net130),
    .B(clknet_1_1__leaf_net355),
    .C(net357),
    .D(net358),
    .Y(net359));
 sky130_fd_sc_hd__nor3b_4 c557 (.A(net353),
    .B(net928),
    .C_N(net932),
    .Y(net360));
 sky130_fd_sc_hd__and4bb_4 c558 (.A_N(net354),
    .B_N(clknet_1_0__leaf_net359),
    .C(clknet_1_1__leaf_net355),
    .D(net224),
    .X(net361));
 sky130_fd_sc_hd__or3b_1 c559 (.A(net918),
    .B(net354),
    .C_N(net944),
    .X(net362));
 sky130_fd_sc_hd__sdfstp_2 c560 (.CLK(clknet_4_3_0_clk),
    .D(net362),
    .SCD(clknet_1_0__leaf_net355),
    .SCE(clknet_1_0__leaf_net245),
    .SET_B(net966),
    .Q(net363));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(clknet_1_0__leaf_net361),
    .A1(net137),
    .A2(net354),
    .A3(net743),
    .S0(clknet_1_0__leaf_net360),
    .S1(net353),
    .X(net364));
 sky130_fd_sc_hd__or3_2 c562 (.A(net363),
    .B(clknet_1_0__leaf_net359),
    .C(net630),
    .X(net365));
 sky130_fd_sc_hd__inv_2 c563 (.A(net579),
    .Y(net366));
 sky130_fd_sc_hd__mux4_2 c564 (.A0(net255),
    .A1(net353),
    .A2(net931),
    .A3(net363),
    .S0(net889),
    .S1(net691),
    .X(net367));
 sky130_fd_sc_hd__nor3_1 c565 (.A(clknet_1_1__leaf_net361),
    .B(net655),
    .C(net692),
    .Y(net368));
 sky130_fd_sc_hd__nor3_1 c566 (.A(clknet_1_1__leaf_net368),
    .B(net362),
    .C(net251),
    .Y(net369));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(net227),
    .A1(net886),
    .A2(clknet_1_0__leaf_net359),
    .A3(net915),
    .S0(net921),
    .S1(net692),
    .X(net370));
 sky130_fd_sc_hd__or3_1 c568 (.A(clknet_1_0__leaf_net368),
    .B(net600),
    .C(clknet_1_1__leaf_net693),
    .X(net371));
 sky130_fd_sc_hd__mux4_4 c569 (.A0(net356),
    .A1(clknet_1_0__leaf_net371),
    .A2(net218),
    .A3(clknet_1_0__leaf_net368),
    .S0(net921),
    .S1(clknet_1_1__leaf_net693),
    .X(net372));
 sky130_fd_sc_hd__mux4_4 c570 (.A0(clknet_1_1__leaf_net371),
    .A1(clknet_1_1__leaf_net365),
    .A2(clknet_1_1__leaf_net368),
    .A3(clknet_1_1__leaf_net372),
    .S0(clknet_1_1__leaf_net220),
    .S1(net692),
    .X(net373));
 sky130_fd_sc_hd__sedfxbp_1 c571 (.CLK(clknet_4_3_0_clk),
    .D(clknet_1_1__leaf_net369),
    .DE(clknet_1_1__leaf_net372),
    .SCD(net972),
    .SCE(clknet_1_0__leaf_net694),
    .Q(net375),
    .Q_N(net374));
 sky130_fd_sc_hd__nand3b_4 c572 (.A_N(net269),
    .B(net153),
    .C(net634),
    .Y(net376));
 sky130_fd_sc_hd__clkbuf_2 c573 (.A(net631),
    .X(net377));
 sky130_fd_sc_hd__or3_2 c574 (.A(net930),
    .B(net272),
    .C(net374),
    .X(net378));
 sky130_fd_sc_hd__sedfxbp_1 c575 (.CLK(clknet_4_12_0_clk),
    .D(net54),
    .DE(net39),
    .SCD(clknet_1_1__leaf_net372),
    .SCE(net890),
    .Q(net380),
    .Q_N(net379));
 sky130_fd_sc_hd__mux4_2 c576 (.A0(net908),
    .A1(net272),
    .A2(net264),
    .A3(net269),
    .S0(net39),
    .S1(clknet_1_0__leaf_net694),
    .X(net381));
 sky130_fd_sc_hd__a2111oi_4 c577 (.A1(net924),
    .A2(clknet_1_1__leaf_net359),
    .B1(net991),
    .C1(net743),
    .D1(net873),
    .Y(net382));
 sky130_fd_sc_hd__and4_2 c578 (.A(clknet_1_0__leaf_net381),
    .B(clknet_1_1__leaf_net161),
    .C(net264),
    .D(clknet_1_1__leaf_net693),
    .X(net858));
 sky130_fd_sc_hd__o2111a_1 c579 (.A1(clknet_1_0__leaf_net382),
    .A2(net224),
    .B1(clknet_1_1__leaf_net161),
    .C1(net376),
    .D1(net914),
    .X(net383));
 sky130_fd_sc_hd__o2111a_2 c580 (.A1(net247),
    .A2(net991),
    .B1(net376),
    .C1(clknet_1_0__leaf_net383),
    .D1(clknet_1_0__leaf_net378),
    .X(net384));
 sky130_fd_sc_hd__nand3_2 c581 (.A(net251),
    .B(net375),
    .C(net923),
    .Y(net385));
 sky130_fd_sc_hd__o2111a_4 c582 (.A1(net264),
    .A2(clknet_1_1__leaf_net361),
    .B1(net239),
    .C1(net914),
    .D1(clknet_1_0__leaf_net383),
    .X(net386));
 sky130_fd_sc_hd__o2111ai_1 c583 (.A1(net385),
    .A2(net887),
    .B1(net891),
    .C1(net908),
    .D1(net615),
    .Y(net387));
 sky130_fd_sc_hd__a2111oi_4 c584 (.A1(clknet_1_1__leaf_net161),
    .A2(clknet_1_0__leaf_net167),
    .B1(net379),
    .C1(net914),
    .D1(net889),
    .Y(net388));
 sky130_fd_sc_hd__sdfbbp_1 c585 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_1__leaf_net372),
    .RESET_B(clknet_1_1__leaf_net382),
    .SCD(clknet_1_1__leaf_net381),
    .SCE(net822),
    .SET_B(clknet_1_1__leaf_net694),
    .Q(net390),
    .Q_N(net389));
 sky130_fd_sc_hd__sdfbbn_2 c586 (.CLK_N(clknet_4_9_0_clk),
    .D(net385),
    .RESET_B(net264),
    .SCD(net39),
    .SCE(clknet_1_1__leaf_net372),
    .SET_B(net890),
    .Q(net392),
    .Q_N(net391));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net890),
    .A1(net389),
    .A2(clknet_1_1__leaf_net167),
    .A3(clknet_1_0__leaf_net383),
    .S0(net615),
    .S1(net637),
    .X(net393));
 sky130_fd_sc_hd__mux4_2 c588 (.A0(net927),
    .A1(net914),
    .A2(net257),
    .A3(net391),
    .S0(net617),
    .S1(clknet_1_0__leaf_net695),
    .X(net832));
 sky130_fd_sc_hd__mux4_4 c589 (.A0(net907),
    .A1(net247),
    .A2(clknet_1_0__leaf_net832),
    .A3(net392),
    .S0(clknet_1_1__leaf_net161),
    .S1(clknet_1_1__leaf_net625),
    .X(net394));
 sky130_fd_sc_hd__a2111oi_2 c590 (.A1(net269),
    .A2(net257),
    .B1(net389),
    .C1(net637),
    .D1(clknet_1_1__leaf_net695),
    .Y(net395));
 sky130_fd_sc_hd__o2111ai_4 c591 (.A1(clknet_1_0__leaf_net395),
    .A2(net914),
    .B1(net907),
    .C1(clknet_1_0__leaf_net832),
    .D1(clknet_1_0__leaf_net695),
    .Y(net396));
 sky130_fd_sc_hd__mux4_2 c592 (.A0(clknet_1_1__leaf_net220),
    .A1(clknet_1_0__leaf_net396),
    .A2(net385),
    .A3(clknet_1_0__leaf_net832),
    .S0(net670),
    .S1(clknet_1_1__leaf_net695),
    .X(net397));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net394),
    .A1(net397),
    .A2(net390),
    .A3(clknet_1_1__leaf_net396),
    .S0(net146),
    .S1(clknet_1_1__leaf_net395),
    .X(net398));
 sky130_fd_sc_hd__buf_8 c594 (.A(clknet_1_0__leaf_net713),
    .X(net399));
 sky130_fd_sc_hd__a2111oi_4 c595 (.A1(net800),
    .A2(clknet_1_1__leaf_net182),
    .B1(net944),
    .C1(net654),
    .D1(net922),
    .Y(net400));
 sky130_fd_sc_hd__buf_12 c596 (.A(clknet_1_1__leaf_net713),
    .X(net401));
 sky130_fd_sc_hd__sedfxtp_4 c597 (.CLK(clknet_4_11_0_clk),
    .D(clknet_1_1__leaf_net245),
    .DE(clknet_1_1__leaf_net399),
    .SCD(clknet_1_1__leaf_net182),
    .SCE(net922),
    .Q(net402));
 sky130_fd_sc_hd__mux4_4 c598 (.A0(net800),
    .A1(net385),
    .A2(clknet_1_1__leaf_net360),
    .A3(clknet_1_1__leaf_net383),
    .S0(net402),
    .S1(net654),
    .X(net403));
 sky130_fd_sc_hd__or3b_2 c599 (.A(clknet_1_0__leaf_net360),
    .B(clknet_1_0__leaf_net399),
    .C_N(net146),
    .X(net404));
 sky130_fd_sc_hd__and3b_1 c600 (.A_N(net380),
    .B(clknet_1_1__leaf_net154),
    .C(net653),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(clknet_1_0__leaf_net404),
    .A1(net908),
    .A2(clknet_1_0__leaf_net858),
    .A3(clknet_1_0__leaf_net399),
    .S0(net653),
    .S1(net816),
    .X(net406));
 sky130_fd_sc_hd__a2111oi_2 c602 (.A1(clknet_1_1__leaf_net399),
    .A2(net402),
    .B1(net887),
    .C1(net377),
    .D1(clknet_1_0__leaf_net677),
    .Y(net407));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net887),
    .A1(net392),
    .A2(net654),
    .A3(net662),
    .S0(net698),
    .S1(net700),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net401),
    .A1(net385),
    .A2(net402),
    .A3(net925),
    .S0(net699),
    .S1(net814),
    .X(net409));
 sky130_fd_sc_hd__mux4_4 c605 (.A0(net409),
    .A1(net375),
    .A2(net249),
    .A3(net377),
    .S0(net303),
    .S1(net816),
    .X(net821));
 sky130_fd_sc_hd__mux4_4 c606 (.A0(clknet_1_1__leaf_net360),
    .A1(net392),
    .A2(clknet_1_0__leaf_net399),
    .A3(net385),
    .S0(clknet_1_1__leaf_net625),
    .S1(net814),
    .X(net410));
 sky130_fd_sc_hd__buf_1 c607 (.A(net715),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net405),
    .A1(clknet_1_0__leaf_net821),
    .A2(net925),
    .A3(net277),
    .S0(net910),
    .S1(net663),
    .X(net412));
 sky130_fd_sc_hd__and3_4 c609 (.A(net411),
    .B(net249),
    .C(net674),
    .X(net413));
 sky130_fd_sc_hd__inv_2 c610 (.A(net875),
    .Y(net414));
 sky130_fd_sc_hd__nand4_4 c611 (.A(net284),
    .B(net249),
    .C(clknet_1_1__leaf_net410),
    .D(net671),
    .Y(net415));
 sky130_fd_sc_hd__inv_6 c612 (.A(net875),
    .Y(net416));
 sky130_fd_sc_hd__mux4_2 c613 (.A0(clknet_1_1__leaf_net378),
    .A1(net277),
    .A2(net411),
    .A3(net413),
    .S0(net416),
    .S1(net402),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net413),
    .A1(clknet_1_1__leaf_net417),
    .A2(clknet_1_1__leaf_net404),
    .A3(net947),
    .S0(net925),
    .S1(net875),
    .X(net418));
 sky130_fd_sc_hd__inv_2 c615 (.A(net716),
    .Y(net825));
 sky130_fd_sc_hd__o2111a_1 c616 (.A1(net91),
    .A2(net99),
    .B1(net791),
    .C1(net96),
    .D1(net312),
    .X(net419));
 sky130_fd_sc_hd__sdfbbn_1 c617 (.CLK_N(clknet_4_14_0_clk),
    .D(net277),
    .RESET_B(net419),
    .SCD(clknet_1_1__leaf_net156),
    .SCE(clknet_1_1__leaf_net182),
    .SET_B(net990),
    .Q(net421),
    .Q_N(net420));
 sky130_fd_sc_hd__o2111a_4 c618 (.A1(clknet_1_1__leaf_net156),
    .A2(net421),
    .B1(net416),
    .C1(net277),
    .D1(clknet_1_1__leaf_net294),
    .X(net422));
 sky130_fd_sc_hd__a2111oi_4 c619 (.A1(net412),
    .A2(net928),
    .B1(clknet_1_0__leaf_net316),
    .C1(net921),
    .D1(net814),
    .Y(net423));
 sky130_fd_sc_hd__a2111oi_2 c620 (.A1(net400),
    .A2(net817),
    .B1(net822),
    .C1(net684),
    .D1(net698),
    .Y(net424));
 sky130_fd_sc_hd__mux4_2 c621 (.A0(clknet_1_1__leaf_net182),
    .A1(net99),
    .A2(net749),
    .A3(net944),
    .S0(net640),
    .S1(net817),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net421),
    .A1(clknet_1_0__leaf_net316),
    .A2(net277),
    .A3(clknet_1_1__leaf_net182),
    .S0(net926),
    .S1(net687),
    .X(net426));
 sky130_fd_sc_hd__o2111a_1 c623 (.A1(clknet_1_1__leaf_net294),
    .A2(clknet_1_0__leaf_net821),
    .B1(net791),
    .C1(clknet_1_1__leaf_net298),
    .D1(net687),
    .X(net427));
 sky130_fd_sc_hd__mux4_2 c624 (.A0(clknet_1_1__leaf_net383),
    .A1(net948),
    .A2(net420),
    .A3(clknet_1_1__leaf_net182),
    .S0(net640),
    .S1(net922),
    .X(net428));
 sky130_fd_sc_hd__a2111o_4 c625 (.A1(net416),
    .A2(net421),
    .B1(net819),
    .C1(net729),
    .D1(clknet_1_1__leaf_net294),
    .X(net429));
 sky130_fd_sc_hd__mux4_2 c626 (.A0(net744),
    .A1(clknet_1_0__leaf_net316),
    .A2(net420),
    .A3(net718),
    .S0(net819),
    .S1(net645),
    .X(net430));
 sky130_fd_sc_hd__mux4_4 c627 (.A0(clknet_1_0__leaf_net298),
    .A1(net926),
    .A2(clknet_1_1__leaf_net156),
    .A3(net958),
    .S0(clknet_1_1__leaf_net425),
    .S1(net920),
    .X(net431));
 sky130_fd_sc_hd__mux4_4 c628 (.A0(clknet_1_0__leaf_net425),
    .A1(clknet_1_1__leaf_net156),
    .A2(net416),
    .A3(net391),
    .S0(net814),
    .S1(net701),
    .X(net432));
 sky130_fd_sc_hd__o2111a_4 c629 (.A1(net946),
    .A2(clknet_1_1__leaf_net182),
    .B1(clknet_1_1__leaf_net832),
    .C1(net822),
    .D1(net818),
    .X(net815));
 sky130_fd_sc_hd__a2111oi_0 c630 (.A1(clknet_1_1__leaf_net182),
    .A2(clknet_1_1__leaf_net815),
    .B1(net865),
    .C1(net850),
    .D1(net920),
    .Y(net433));
 sky130_fd_sc_hd__mux4_2 c631 (.A0(net925),
    .A1(clknet_1_0__leaf_net815),
    .A2(clknet_1_1__leaf_net156),
    .A3(clknet_1_1__leaf_net425),
    .S0(net684),
    .S1(net701),
    .X(net434));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net390),
    .A1(clknet_1_0__leaf_net425),
    .A2(clknet_1_1__leaf_net815),
    .A3(net416),
    .S0(net670),
    .S1(net702),
    .X(net435));
 sky130_fd_sc_hd__mux4_4 c633 (.A0(clknet_1_1__leaf_net435),
    .A1(net313),
    .A2(clknet_1_0__leaf_net316),
    .A3(clknet_1_0__leaf_net815),
    .S0(net684),
    .S1(net702),
    .X(net436));
 sky130_fd_sc_hd__mux4_4 c634 (.A0(clknet_1_0__leaf_net435),
    .A1(clknet_1_1__leaf_net821),
    .A2(net791),
    .A3(clknet_1_1__leaf_net424),
    .S0(net817),
    .S1(net702),
    .X(net824));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net433),
    .A1(clknet_1_1__leaf_net298),
    .A2(clknet_1_1__leaf_net435),
    .A3(net850),
    .S0(net920),
    .S1(net702),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(clknet_1_0__leaf_net424),
    .A1(clknet_1_0__leaf_net435),
    .A2(net925),
    .A3(net645),
    .S0(net649),
    .S1(net702),
    .X(net823));
 sky130_fd_sc_hd__mux4_4 c637 (.A0(net99),
    .A1(net841),
    .A2(net420),
    .A3(clknet_1_0__leaf_net815),
    .S0(net649),
    .S1(net702),
    .X(net438));
 sky130_fd_sc_hd__or2b_1 c660 (.A(net915),
    .B_N(net586),
    .X(net439));
 sky130_fd_sc_hd__nor2_2 c661 (.A(net217),
    .B(net343),
    .Y(net440));
 sky130_fd_sc_hd__nor2_1 c662 (.A(net439),
    .B(net648),
    .Y(net441));
 sky130_fd_sc_hd__or3_2 c663 (.A(net441),
    .B(net909),
    .C(net690),
    .X(net442));
 sky130_fd_sc_hd__nor2b_1 c664 (.A(net440),
    .B_N(net442),
    .Y(net443));
 sky130_fd_sc_hd__nor2b_1 c665 (.A(net350),
    .B_N(net343),
    .Y(net444));
 sky130_fd_sc_hd__and2_1 c666 (.A(net439),
    .B(net586),
    .X(net445));
 sky130_fd_sc_hd__or3b_1 c667 (.A(net444),
    .B(net442),
    .C_N(net440),
    .X(net446));
 sky130_fd_sc_hd__or3b_2 c668 (.A(net343),
    .B(net439),
    .C_N(net444),
    .X(net447));
 sky130_fd_sc_hd__buf_6 c669 (.A(net596),
    .X(net448));
 sky130_fd_sc_hd__nand4b_4 c670 (.A_N(net440),
    .B(net927),
    .C(net447),
    .D(net690),
    .Y(net449));
 sky130_fd_sc_hd__sedfxtp_4 c671 (.CLK(clknet_4_2_0_clk),
    .D(net442),
    .DE(clknet_1_0__leaf_net337),
    .SCD(net905),
    .SCE(net448),
    .Q(net450));
 sky130_fd_sc_hd__nor3_1 c672 (.A(net448),
    .B(net445),
    .C(net905),
    .Y(net451));
 sky130_fd_sc_hd__mux4_2 c673 (.A0(net446),
    .A1(net440),
    .A2(net905),
    .A3(net109),
    .S0(net586),
    .S1(net688),
    .X(net452));
 sky130_fd_sc_hd__nand3_1 c674 (.A(net113),
    .B(net349),
    .C(net443),
    .Y(net453));
 sky130_fd_sc_hd__nor3_1 c675 (.A(net218),
    .B(net440),
    .C(net442),
    .Y(net454));
 sky130_fd_sc_hd__and4b_1 c676 (.A_N(net453),
    .B(net454),
    .C(net442),
    .D(net445),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_2 c677 (.A(net596),
    .X(net456));
 sky130_fd_sc_hd__nor3_2 c678 (.A(net455),
    .B(net440),
    .C(net454),
    .Y(net457));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net451),
    .A1(net113),
    .A2(net456),
    .A3(net915),
    .S0(net109),
    .S1(net689),
    .X(net458));
 sky130_fd_sc_hd__sedfxtp_2 c680 (.CLK(clknet_4_2_0_clk),
    .D(net443),
    .DE(net457),
    .SCD(net455),
    .SCE(net458),
    .Q(net459));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net458),
    .A1(net453),
    .A2(net441),
    .A3(net439),
    .S0(net343),
    .S1(net459),
    .X(net460));
 sky130_fd_sc_hd__a2111oi_2 c682 (.A1(net450),
    .A2(net926),
    .B1(net905),
    .C1(net927),
    .D1(net668),
    .Y(net461));
 sky130_fd_sc_hd__sdfbbp_1 c683 (.CLK(clknet_4_2_0_clk),
    .D(net366),
    .RESET_B(net457),
    .SCD(net456),
    .SCE(net445),
    .SET_B(net969),
    .Q(net463),
    .Q_N(net462));
 sky130_fd_sc_hd__sdfbbn_1 c684 (.CLK_N(clknet_4_2_0_clk),
    .D(net459),
    .RESET_B(net990),
    .SCD(net905),
    .SCE(net457),
    .SET_B(net597),
    .Q(net465),
    .Q_N(net464));
 sky130_fd_sc_hd__sdfrbp_1 c685 (.CLK(clknet_4_2_0_clk),
    .D(net125),
    .RESET_B(net962),
    .SCD(net366),
    .SCE(net464),
    .Q(net467),
    .Q_N(net466));
 sky130_fd_sc_hd__o2111ai_4 c686 (.A1(net456),
    .A2(net465),
    .B1(net239),
    .C1(net926),
    .D1(net450),
    .Y(net468));
 sky130_fd_sc_hd__sdfbbn_2 c687 (.CLK_N(clknet_4_2_0_clk),
    .D(net445),
    .RESET_B(net457),
    .SCD(net459),
    .SCE(net363),
    .SET_B(net921),
    .Q(net470),
    .Q_N(net469));
 sky130_fd_sc_hd__mux4_2 c688 (.A0(net463),
    .A1(net465),
    .A2(net743),
    .A3(net467),
    .S0(net905),
    .S1(net468),
    .X(net471));
 sky130_fd_sc_hd__nor3_2 c689 (.A(net109),
    .B(net468),
    .C(net239),
    .Y(net472));
 sky130_fd_sc_hd__mux4_4 c690 (.A0(net462),
    .A1(clknet_1_0__leaf_net369),
    .A2(net471),
    .A3(net470),
    .S0(net256),
    .S1(net597),
    .X(net473));
 sky130_fd_sc_hd__inv_2 c691 (.A(net647),
    .Y(net474));
 sky130_fd_sc_hd__or4_1 c692 (.A(net457),
    .B(net463),
    .C(net470),
    .D(net456),
    .X(net475));
 sky130_fd_sc_hd__nand3_4 c693 (.A(net363),
    .B(net461),
    .C(net464),
    .Y(net476));
 sky130_fd_sc_hd__a2111oi_1 c694 (.A1(clknet_1_0__leaf_net355),
    .A2(net915),
    .B1(net470),
    .C1(net356),
    .D1(net891),
    .Y(net477));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net357),
    .A1(net471),
    .A2(net472),
    .A3(net466),
    .S0(net474),
    .S1(net356),
    .X(net478));
 sky130_fd_sc_hd__o2111ai_4 c696 (.A1(net257),
    .A2(net356),
    .B1(net918),
    .C1(net469),
    .D1(net643),
    .Y(net479));
 sky130_fd_sc_hd__inv_1 c697 (.A(net647),
    .Y(net480));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net467),
    .A1(net462),
    .A2(net915),
    .A3(net465),
    .S0(net480),
    .S1(net643),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net356),
    .A1(net905),
    .A2(net480),
    .A3(net481),
    .S0(net472),
    .S1(net331),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net470),
    .A1(net33),
    .A2(net480),
    .A3(net331),
    .S0(net452),
    .S1(net468),
    .X(net483));
 sky130_fd_sc_hd__mux4_2 c701 (.A0(net481),
    .A1(net480),
    .A2(net466),
    .A3(net905),
    .S0(net634),
    .S1(clknet_1_0__leaf_net693),
    .X(net484));
 sky130_fd_sc_hd__mux4_4 c702 (.A0(net479),
    .A1(net481),
    .A2(net456),
    .A3(net480),
    .S0(net476),
    .S1(clknet_1_0__leaf_net484),
    .X(net485));
 sky130_fd_sc_hd__mux4_2 c703 (.A0(net485),
    .A1(net480),
    .A2(net481),
    .A3(clknet_1_0__leaf_net372),
    .S0(net729),
    .S1(net469),
    .X(net486));
 sky130_fd_sc_hd__mux4_4 c704 (.A0(net890),
    .A1(net392),
    .A2(clknet_1_0__leaf_net477),
    .A3(net914),
    .S0(net614),
    .S1(clknet_1_0__leaf_net693),
    .X(net487));
 sky130_fd_sc_hd__and3b_1 c705 (.A_N(clknet_1_0__leaf_net484),
    .B(net146),
    .C(net672),
    .X(net488));
 sky130_fd_sc_hd__mux4_4 c706 (.A0(net239),
    .A1(net991),
    .A2(clknet_1_0__leaf_net372),
    .A3(clknet_1_0__leaf_net477),
    .S0(net479),
    .S1(net391),
    .X(net489));
 sky130_fd_sc_hd__sdfbbp_1 c707 (.CLK(clknet_4_8_0_clk),
    .D(net993),
    .RESET_B(net39),
    .SCD(net452),
    .SCE(clknet_1_0__leaf_net372),
    .SET_B(clknet_1_0__leaf_net231),
    .Q(net491),
    .Q_N(net490));
 sky130_fd_sc_hd__a2111oi_2 c708 (.A1(net923),
    .A2(net479),
    .B1(net918),
    .C1(net145),
    .D1(net671),
    .Y(net492));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net473),
    .A1(net491),
    .A2(net146),
    .A3(net452),
    .S0(net376),
    .S1(net671),
    .X(net493));
 sky130_fd_sc_hd__sdfbbn_1 c710 (.CLK_N(clknet_4_8_0_clk),
    .D(net452),
    .RESET_B(net749),
    .SCD(clknet_1_0__leaf_net477),
    .SCE(net648),
    .SET_B(net671),
    .Q(net495),
    .Q_N(net494));
 sky130_fd_sc_hd__a2111oi_1 c711 (.A1(net376),
    .A2(net479),
    .B1(net476),
    .C1(net668),
    .D1(net703),
    .Y(net496));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net979),
    .A1(net376),
    .A2(net890),
    .A3(net906),
    .S0(net672),
    .S1(net703),
    .X(net497));
 sky130_fd_sc_hd__o2111a_4 c713 (.A1(net495),
    .A2(net890),
    .B1(net490),
    .C1(clknet_1_1__leaf_net484),
    .D1(clknet_1_0__leaf_net693),
    .X(net498));
 sky130_fd_sc_hd__mux4_4 c714 (.A0(net471),
    .A1(net488),
    .A2(net887),
    .A3(net479),
    .S0(net896),
    .S1(net671),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net498),
    .A1(net494),
    .A2(net238),
    .A3(net648),
    .S0(net672),
    .S1(net704),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net491),
    .A1(net923),
    .A2(net890),
    .A3(net39),
    .S0(net671),
    .S1(net697),
    .X(net501));
 sky130_fd_sc_hd__sdfbbn_1 c717 (.CLK_N(clknet_4_8_0_clk),
    .D(net452),
    .RESET_B(net471),
    .SCD(net973),
    .SCE(net703),
    .SET_B(net704),
    .Q(net503),
    .Q_N(net502));
 sky130_fd_sc_hd__sdfbbp_1 c718 (.CLK(clknet_4_8_0_clk),
    .D(net890),
    .RESET_B(net503),
    .SCD(net903),
    .SCE(net452),
    .SET_B(net965),
    .Q(net505),
    .Q_N(net504));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net744),
    .A1(net492),
    .A2(net472),
    .A3(clknet_1_0__leaf_net231),
    .S0(net479),
    .S1(net923),
    .X(net506));
 sky130_fd_sc_hd__mux4_4 c720 (.A0(net472),
    .A1(net505),
    .A2(net491),
    .A3(net470),
    .S0(net624),
    .S1(net641),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net501),
    .A1(net890),
    .A2(net472),
    .A3(net744),
    .S0(net504),
    .S1(net641),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net480),
    .A1(net903),
    .A2(net501),
    .A3(net624),
    .S0(net703),
    .S1(net706),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net497),
    .A1(net502),
    .A2(net490),
    .A3(net902),
    .S0(net914),
    .S1(net706),
    .X(net510));
 sky130_fd_sc_hd__mux4_4 c724 (.A0(clknet_1_0__leaf_net372),
    .A1(net902),
    .A2(net614),
    .A3(net647),
    .S0(net672),
    .S1(net705),
    .X(net511));
 sky130_fd_sc_hd__sdfrbp_1 c725 (.CLK(clknet_4_8_0_clk),
    .D(net472),
    .RESET_B(net890),
    .SCD(net624),
    .SCE(net709),
    .Q(net513),
    .Q_N(net512));
 sky130_fd_sc_hd__o2111a_1 c726 (.A1(net413),
    .A2(net928),
    .B1(net6),
    .C1(net918),
    .D1(net391),
    .X(net514));
 sky130_fd_sc_hd__o2111ai_1 c727 (.A1(net514),
    .A2(net905),
    .B1(net513),
    .C1(clknet_1_0__leaf_net477),
    .D1(net729),
    .Y(net515));
 sky130_fd_sc_hd__mux4_4 c728 (.A0(net402),
    .A1(net749),
    .A2(net743),
    .A3(net238),
    .S0(net33),
    .S1(net708),
    .X(net516));
 sky130_fd_sc_hd__mux4_2 c729 (.A0(net474),
    .A1(net176),
    .A2(net449),
    .A3(net745),
    .S0(net672),
    .S1(net921),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net896),
    .A1(net304),
    .A2(net413),
    .A3(net474),
    .S0(net887),
    .S1(net671),
    .X(net518));
 sky130_fd_sc_hd__o2111ai_4 c731 (.A1(net476),
    .A2(net402),
    .B1(net413),
    .C1(net928),
    .D1(net708),
    .Y(net519));
 sky130_fd_sc_hd__o2111ai_4 c732 (.A1(net517),
    .A2(net146),
    .B1(net238),
    .C1(net469),
    .D1(net674),
    .Y(net520));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net449),
    .A1(net238),
    .A2(net256),
    .A3(net519),
    .S0(net413),
    .S1(net708),
    .X(net521));
 sky130_fd_sc_hd__o2111ai_1 c734 (.A1(net225),
    .A2(net33),
    .B1(net391),
    .C1(net512),
    .D1(net672),
    .Y(net522));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net519),
    .A1(net303),
    .A2(net922),
    .A3(net672),
    .S0(net674),
    .S1(net921),
    .X(net523));
 sky130_fd_sc_hd__mux4_4 c736 (.A0(net523),
    .A1(net303),
    .A2(net887),
    .A3(net469),
    .S0(net672),
    .S1(net707),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net520),
    .A1(net519),
    .A2(net599),
    .A3(net671),
    .S0(net691),
    .S1(net707),
    .X(net525));
 sky130_fd_sc_hd__mux4_2 c738 (.A0(net525),
    .A1(net519),
    .A2(net905),
    .A3(net943),
    .S0(net636),
    .S1(net671),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net516),
    .A1(net513),
    .A2(net176),
    .A3(net519),
    .S0(net672),
    .S1(net707),
    .X(net527));
 sky130_fd_sc_hd__mux4_4 c740 (.A0(net522),
    .A1(net520),
    .A2(net33),
    .A3(net238),
    .S0(net674),
    .S1(net709),
    .X(net528));
 sky130_fd_sc_hd__mux4_4 c741 (.A0(net257),
    .A1(net519),
    .A2(net523),
    .A3(net402),
    .S0(net526),
    .S1(net672),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net528),
    .A1(net470),
    .A2(net527),
    .A3(net519),
    .S0(net525),
    .S1(net709),
    .X(net530));
 sky130_fd_sc_hd__mux4_4 c743 (.A0(net238),
    .A1(net530),
    .A2(net527),
    .A3(net520),
    .S0(net256),
    .S1(net523),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net530),
    .A1(net520),
    .A2(net413),
    .A3(net743),
    .S0(net634),
    .S1(net696),
    .X(net532));
 sky130_fd_sc_hd__mux4_4 c745 (.A0(net527),
    .A1(net402),
    .A2(net526),
    .A3(net525),
    .S0(net710),
    .S1(net711),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net887),
    .A1(net33),
    .A2(net469),
    .A3(net646),
    .S0(net710),
    .S1(net711),
    .X(net534));
 sky130_fd_sc_hd__mux4_2 c747 (.A0(net928),
    .A1(net413),
    .A2(net28),
    .A3(net256),
    .S0(clknet_1_0__leaf_net627),
    .S1(net646),
    .X(net535));
 sky130_fd_sc_hd__mux4_2 c748 (.A0(clknet_1_1__leaf_net417),
    .A1(net526),
    .A2(clknet_1_1__leaf_net477),
    .A3(net599),
    .S0(net696),
    .S1(net709),
    .X(net536));
 sky130_fd_sc_hd__mux4_2 c749 (.A0(net392),
    .A1(net914),
    .A2(clknet_1_1__leaf_net477),
    .A3(clknet_1_1__leaf_net417),
    .S0(net920),
    .S1(net709),
    .X(net537));
 sky130_fd_sc_hd__mux4_4 c750 (.A0(net535),
    .A1(net928),
    .A2(net943),
    .A3(net729),
    .S0(net921),
    .S1(net920),
    .X(net538));
 sky130_fd_sc_hd__mux4_4 c751 (.A0(net928),
    .A1(net512),
    .A2(net526),
    .A3(net650),
    .S0(net920),
    .S1(net711),
    .X(net539));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net513),
    .A1(clknet_1_0__leaf_net231),
    .A2(net526),
    .A3(net6),
    .S0(clknet_1_0__leaf_net477),
    .S1(net920),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net313),
    .A1(net943),
    .A2(net650),
    .A3(net922),
    .S0(net920),
    .S1(net711),
    .X(net541));
 sky130_fd_sc_hd__mux4_4 c754 (.A0(clknet_1_1__leaf_net477),
    .A1(net521),
    .A2(net313),
    .A3(net526),
    .S0(net921),
    .S1(net709),
    .X(net542));
 sky130_fd_sc_hd__mux4_4 c755 (.A0(net914),
    .A1(clknet_1_0__leaf_net417),
    .A2(net512),
    .A3(clknet_1_1__leaf_net477),
    .S0(net640),
    .S1(net711),
    .X(net543));
 sky130_fd_sc_hd__mux4_4 c756 (.A0(net96),
    .A1(clknet_1_1__leaf_net417),
    .A2(net691),
    .A3(net697),
    .S0(net709),
    .S1(net711),
    .X(net544));
 sky130_fd_sc_hd__mux4_4 c757 (.A0(net526),
    .A1(net749),
    .A2(net312),
    .A3(net641),
    .S0(net668),
    .S1(net711),
    .X(net545));
 sky130_fd_sc_hd__mux4_2 c758 (.A0(clknet_1_0__leaf_net417),
    .A1(clknet_1_1__leaf_net477),
    .A2(net312),
    .A3(net641),
    .S0(net642),
    .S1(net920),
    .X(net546));
 sky130_fd_sc_hd__mux4_2 c759 (.A0(net526),
    .A1(clknet_1_0__leaf_net417),
    .A2(net914),
    .A3(net312),
    .S0(net642),
    .S1(clknet_1_0__leaf_net712),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net313),
    .A1(net541),
    .A2(clknet_1_1__leaf_net477),
    .A3(net526),
    .S0(net650),
    .S1(net711),
    .X(net548));
 sky130_fd_sc_hd__mux4_2 c761 (.A0(clknet_1_0__leaf_net231),
    .A1(clknet_1_0__leaf_net417),
    .A2(clknet_1_1__leaf_net627),
    .A3(net650),
    .S0(net920),
    .S1(clknet_1_1__leaf_net712),
    .X(net549));
 sky130_fd_sc_hd__mux4_2 c762 (.A0(net538),
    .A1(net613),
    .A2(net636),
    .A3(net921),
    .S0(net711),
    .S1(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__mux4_1 merge763 (.A0(net53),
    .A1(net35),
    .A2(net50),
    .A3(net56),
    .S0(net58),
    .S1(net620),
    .X(net550));
 sky130_fd_sc_hd__mux4_1 merge764 (.A0(net211),
    .A1(net214),
    .A2(net885),
    .A3(clknet_1_0__leaf_net228),
    .S0(net216),
    .S1(clknet_1_1__leaf_net229),
    .X(net551));
 sky130_fd_sc_hd__mux4_1 merge765 (.A0(net177),
    .A1(net945),
    .A2(net910),
    .A3(net238),
    .S0(clknet_1_0__leaf_net298),
    .S1(clknet_1_0__leaf_net677),
    .X(net552));
 sky130_fd_sc_hd__o2111a_1 merge766 (.A1(net863),
    .A2(net55),
    .B1(net767),
    .C1(net53),
    .D1(net603),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 merge767 (.A0(net152),
    .A1(clknet_1_0__leaf_net157),
    .A2(net886),
    .A3(clknet_1_0__leaf_net161),
    .S0(clknet_1_0__leaf_net156),
    .S1(net132),
    .X(net554));
 sky130_fd_sc_hd__mux4_4 merge768 (.A0(net747),
    .A1(net886),
    .A2(net129),
    .A3(net45),
    .S0(net136),
    .S1(net585),
    .X(net555));
 sky130_fd_sc_hd__a2111oi_2 merge769 (.A1(net732),
    .A2(net243),
    .B1(clknet_1_1__leaf_net151),
    .C1(net892),
    .D1(net134),
    .Y(net556));
 sky130_fd_sc_hd__mux4_4 merge770 (.A0(net447),
    .A1(net446),
    .A2(net125),
    .A3(net451),
    .S0(net448),
    .S1(clknet_1_0__leaf_net231),
    .X(net557));
 sky130_fd_sc_hd__mux4_4 merge771 (.A0(net915),
    .A1(clknet_1_0__leaf_net231),
    .A2(net330),
    .A3(net332),
    .S0(net334),
    .S1(clknet_1_1__leaf_net657),
    .X(net558));
 sky130_fd_sc_hd__mux4_2 merge772 (.A0(net236),
    .A1(clknet_1_0__leaf_net245),
    .A2(net239),
    .A3(net352),
    .S0(net918),
    .S1(net655),
    .X(net559));
 sky130_fd_sc_hd__mux4_4 merge773 (.A0(net464),
    .A1(clknet_1_0__leaf_net231),
    .A2(net450),
    .A3(net137),
    .S0(net239),
    .S1(net992),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 merge774 (.A0(clknet_1_1__leaf_net165),
    .A1(net886),
    .A2(net250),
    .A3(net762),
    .S0(net883),
    .S1(clknet_1_0__leaf_net156),
    .X(net561));
 sky130_fd_sc_hd__mux4_4 merge775 (.A0(net177),
    .A1(clknet_1_0__leaf_net410),
    .A2(net416),
    .A3(net374),
    .S0(clknet_1_1__leaf_net245),
    .S1(net670),
    .X(net562));
 sky130_fd_sc_hd__a2111o_1 merge776 (.A1(net58),
    .A2(net56),
    .B1(net725),
    .C1(net52),
    .D1(net63),
    .X(net563));
 sky130_fd_sc_hd__mux4_4 merge777 (.A0(clknet_1_1__leaf_net159),
    .A1(clknet_1_0__leaf_net161),
    .A2(net265),
    .A3(net162),
    .S0(net260),
    .S1(net638),
    .X(net564));
 sky130_fd_sc_hd__a2111oi_2 merge778 (.A1(clknet_1_1__leaf_net228),
    .A2(net889),
    .B1(net340),
    .C1(net226),
    .D1(net667),
    .Y(net565));
 sky130_fd_sc_hd__mux4_2 merge779 (.A0(net352),
    .A1(net250),
    .A2(net966),
    .A3(clknet_1_0__leaf_net365),
    .S0(net243),
    .S1(net921),
    .X(net566));
 sky130_fd_sc_hd__mux4_1 merge780 (.A0(net88),
    .A1(net95),
    .A2(net55),
    .A3(net9),
    .S0(net784),
    .S1(net78),
    .X(net567));
 sky130_fd_sc_hd__mux4_2 merge781 (.A0(net884),
    .A1(clknet_1_1__leaf_net231),
    .A2(net908),
    .A3(net162),
    .S0(net960),
    .S1(clknet_1_0__leaf_net361),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(net414),
    .A1(net415),
    .A2(net177),
    .A3(clknet_1_0__leaf_net305),
    .S0(clknet_1_1__leaf_net383),
    .S1(clknet_1_1__leaf_net832),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(net268),
    .A1(net261),
    .A2(net236),
    .A3(net37),
    .S0(net884),
    .S1(net644),
    .X(net570));
 sky130_fd_sc_hd__a2111o_1 merge784 (.A1(net243),
    .A2(net240),
    .B1(clknet_1_1__leaf_net231),
    .C1(net242),
    .D1(net236),
    .X(net571));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net66),
    .A1(net893),
    .A2(clknet_1_0__leaf_net245),
    .A3(net263),
    .S0(net884),
    .S1(net617),
    .X(net572));
 sky130_fd_sc_hd__or2_1 merge786 (.A(net168),
    .B(net171),
    .X(net573));
 sky130_fd_sc_hd__nor2_1 merge787 (.A(net475),
    .B(net478),
    .Y(net574));
 sky130_fd_sc_hd__nor2_1 merge788 (.A(net422),
    .B(net426),
    .Y(net575));
 sky130_fd_sc_hd__or2b_4 merge789 (.A(net407),
    .B_N(net418),
    .X(net576));
 sky130_fd_sc_hd__and2_1 merge790 (.A(net384),
    .B(net387),
    .X(net577));
 sky130_fd_sc_hd__or2b_1 merge791 (.A(net43),
    .B_N(net44),
    .X(net578));
 sky130_fd_sc_hd__dfrbp_2 merge792 (.CLK(clknet_4_3_0_clk),
    .D(net559),
    .RESET_B(net566),
    .Q(net580),
    .Q_N(net579));
 sky130_fd_sc_hd__dfrbp_1 merge793 (.CLK(clknet_4_7_0_clk),
    .D(net189),
    .RESET_B(net175),
    .Q(net582),
    .Q_N(net581));
 sky130_fd_sc_hd__nor2b_2 merge794 (.A(net536),
    .B_N(net537),
    .Y(net583));
 sky130_fd_sc_hd__nor2b_4 merge795 (.A(net315),
    .B_N(net326),
    .Y(net584));
 sky130_fd_sc_hd__dfrtn_1 merge796 (.CLK_N(clknet_4_1_0_clk),
    .D(net122),
    .RESET_B(net111),
    .Q(net585));
 sky130_fd_sc_hd__dfrtp_2 merge797 (.CLK(clknet_4_0_0_clk),
    .D(net551),
    .RESET_B(net234),
    .Q(net586));
 sky130_fd_sc_hd__and2b_1 merge798 (.A_N(net84),
    .B(net85),
    .X(net587));
 sky130_fd_sc_hd__dfrtp_1 merge799 (.CLK(clknet_4_1_0_clk),
    .D(net338),
    .Q(net341));
 sky130_fd_sc_hd__and2b_1 merge800 (.A_N(net200),
    .B(net203),
    .X(net589));
 sky130_fd_sc_hd__and2_1 merge801 (.A(net102),
    .B(net89),
    .X(net590));
 sky130_fd_sc_hd__dfrtp_1 merge802 (.CLK(clknet_4_12_0_clk),
    .D(net290),
    .RESET_B(net300),
    .Q(net591));
 sky130_fd_sc_hd__or2_1 merge803 (.A(net489),
    .B(net509),
    .X(net592));
 sky130_fd_sc_hd__dfsbp_2 merge804 (.CLK(clknet_4_6_0_clk),
    .D(net266),
    .SET_B(net561),
    .Q(net594),
    .Q_N(net593));
 sky130_fd_sc_hd__and2b_1 merge805 (.A_N(net59),
    .B(net550),
    .X(net595));
 sky130_fd_sc_hd__dfsbp_1 merge806 (.CLK(clknet_4_2_0_clk),
    .D(net460),
    .SET_B(net557),
    .Q(net597),
    .Q_N(net596));
 sky130_fd_sc_hd__and2_0 merge807 (.A(net148),
    .B(net149),
    .X(net598));
 sky130_fd_sc_hd__dfstp_1 merge808 (.CLK(clknet_4_9_0_clk),
    .D(net515),
    .SET_B(net518),
    .Q(net599));
 sky130_fd_sc_hd__dfstp_1 merge809 (.CLK(clknet_4_1_0_clk),
    .D(net252),
    .SET_B(net254),
    .Q(net600));
 sky130_fd_sc_hd__nor2b_4 merge810 (.A(net486),
    .B_N(net483),
    .Y(net601));
 sky130_fd_sc_hd__and2_4 merge811 (.A(net329),
    .B(net438),
    .X(net602));
 sky130_fd_sc_hd__dfstp_2 merge812 (.CLK(clknet_4_5_0_clk),
    .D(net563),
    .SET_B(net62),
    .Q(net603));
 sky130_fd_sc_hd__nand2b_1 merge813 (.A_N(net98),
    .B(net567),
    .Y(net604));
 sky130_fd_sc_hd__dlrbn_1 merge814 (.D(net555),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net147),
    .Q(net606),
    .Q_N(net605));
 sky130_fd_sc_hd__or2b_2 merge815 (.A(net427),
    .B_N(net428),
    .X(net607));
 sky130_fd_sc_hd__dlrbn_1 merge816 (.D(net553),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net80),
    .Q(net609),
    .Q_N(net608));
 sky130_fd_sc_hd__dlrbp_1 merge817 (.D(net196),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net584),
    .Q(net610),
    .Q_N(net840));
 sky130_fd_sc_hd__nand2b_1 merge818 (.A_N(net204),
    .B(net208),
    .Y(net611));
 sky130_fd_sc_hd__and2_1 merge819 (.A(net510),
    .B(net549),
    .X(net612));
 sky130_fd_sc_hd__dlrbp_1 merge820 (.D(net482),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net612),
    .Q(net614),
    .Q_N(net613));
 sky130_fd_sc_hd__dlrtn_2 merge821 (.D(net577),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net347),
    .Q(net615));
 sky130_fd_sc_hd__dlrtn_2 merge822 (.D(net571),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net556),
    .Q(net616));
 sky130_fd_sc_hd__dlrtn_1 merge823 (.D(net345),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net259),
    .Q(net617));
 sky130_fd_sc_hd__dlrtp_2 merge824 (.D(net310),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net327),
    .Q(net834));
 sky130_fd_sc_hd__and2_1 merge825 (.A(net529),
    .B(net524),
    .X(net618));
 sky130_fd_sc_hd__and2_2 merge826 (.A(net544),
    .B(net548),
    .X(net619));
 sky130_fd_sc_hd__dlrtp_2 merge827 (.D(net590),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net595),
    .Q(net620));
 sky130_fd_sc_hd__dlrtp_2 merge828 (.D(net587),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net604),
    .Q(net621));
 sky130_fd_sc_hd__edfxbp_1 merge829 (.CLK(clknet_4_5_0_clk),
    .D(net564),
    .DE(net554),
    .Q(net623),
    .Q_N(net622));
 sky130_fd_sc_hd__edfxtp_1 merge830 (.CLK(clknet_4_8_0_clk),
    .D(net592),
    .DE(net506),
    .Q(net624));
 sky130_fd_sc_hd__sdlclkp_1 merge831 (.CLK(clknet_4_6_0_clk),
    .GATE(net598),
    .SCE(net170),
    .GCLK(net625));
 sky130_fd_sc_hd__sdlclkp_2 merge832 (.CLK(clknet_4_4_0_clk),
    .SCE(net578),
    .GCLK(net46));
 sky130_fd_sc_hd__sdlclkp_4 merge833 (.CLK(clknet_4_10_0_clk),
    .GATE(net534),
    .SCE(net547),
    .GCLK(net627));
 sky130_fd_sc_hd__nand2_2 merge834 (.A(net431),
    .B(net432),
    .Y(net628));
 sky130_fd_sc_hd__dfrbp_1 merge835 (.CLK(clknet_4_6_0_clk),
    .D(net258),
    .RESET_B(net572),
    .Q(net630),
    .Q_N(net629));
 sky130_fd_sc_hd__dfrbp_2 merge836 (.CLK(clknet_4_6_0_clk),
    .D(net570),
    .RESET_B(net568),
    .Q(net632),
    .Q_N(net631));
 sky130_fd_sc_hd__dfrtn_1 merge837 (.CLK_N(clknet_4_15_0_clk),
    .D(net325),
    .RESET_B(net209),
    .Q(net830));
 sky130_fd_sc_hd__or2b_1 merge838 (.A(net539),
    .B_N(net546),
    .X(net633));
 sky130_fd_sc_hd__dfrtp_4 merge839 (.CLK(clknet_4_11_0_clk),
    .D(net576),
    .RESET_B(net569),
    .Q(net875));
 sky130_fd_sc_hd__dfrtp_4 merge840 (.CLK(clknet_4_3_0_clk),
    .D(net351),
    .RESET_B(net601),
    .Q(net634));
 sky130_fd_sc_hd__dfrtp_2 merge841 (.CLK(clknet_4_13_0_clk),
    .D(net210),
    .RESET_B(net589),
    .Q(net635));
 sky130_fd_sc_hd__dfsbp_1 merge842 (.CLK(clknet_4_9_0_clk),
    .D(net386),
    .SET_B(net618),
    .Q(net637),
    .Q_N(net636));
 sky130_fd_sc_hd__dfsbp_1 merge843 (.CLK(clknet_4_14_0_clk),
    .D(net628),
    .SET_B(net607),
    .Q(net869),
    .Q_N(net865));
 sky130_fd_sc_hd__dfstp_2 merge844 (.CLK(clknet_4_5_0_clk),
    .D(net185),
    .SET_B(net160),
    .Q(net638));
 sky130_fd_sc_hd__or2b_2 merge845 (.A(net540),
    .B_N(net543),
    .X(net639));
 sky130_fd_sc_hd__dfstp_2 merge846 (.CLK(clknet_4_11_0_clk),
    .D(net542),
    .SET_B(net575),
    .Q(net640));
 sky130_fd_sc_hd__dfstp_1 merge847 (.CLK(clknet_4_10_0_clk),
    .D(net500),
    .SET_B(net639),
    .Q(net641));
 sky130_fd_sc_hd__dlrbn_1 merge848 (.D(net319),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net602),
    .Q(net833),
    .Q_N(net820));
 sky130_fd_sc_hd__dlrbn_1 merge849 (.D(net574),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net633),
    .Q(net643),
    .Q_N(net642));
 sky130_fd_sc_hd__dlrbp_2 merge850 (.D(net169),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net190),
    .Q(net644),
    .Q_N(net839));
 sky130_fd_sc_hd__dlrbp_1 merge851 (.D(net533),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net429),
    .Q(net646),
    .Q_N(net645));
 sky130_fd_sc_hd__dlrtn_1 merge852 (.D(net560),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net487),
    .Q(net647));
 sky130_fd_sc_hd__dlrtn_2 merge853 (.D(net611),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net186),
    .Q(net847));
 sky130_fd_sc_hd__dlrtn_1 merge854 (.D(net348),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net388),
    .Q(net648));
 sky130_fd_sc_hd__dlrtp_4 merge855 (.D(net565),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net437),
    .Q(net649));
 sky130_fd_sc_hd__dlrtp_4 merge856 (.D(net188),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net573),
    .Q(net846));
 sky130_fd_sc_hd__dlrtp_1 merge857 (.D(net619),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net583),
    .Q(net650));
 sky130_fd_sc_hd__edfxbp_1 merge858 (.CLK(clknet_4_13_0_clk),
    .D(net198),
    .DE(net205),
    .Q(net651),
    .Q_N(net842));
 sky130_fd_sc_hd__edfxtp_1 merge859 (.CLK(clknet_4_14_0_clk),
    .D(net436),
    .DE(net423),
    .Q(net817));
 sky130_fd_sc_hd__dfxbp_2 s860 (.CLK(clknet_4_5_0_clk),
    .D(net77),
    .Q(net848),
    .Q_N(net652));
 sky130_fd_sc_hd__dfxbp_2 s861 (.CLK(clknet_4_7_0_clk),
    .D(net82),
    .Q(net654),
    .Q_N(net653));
 sky130_fd_sc_hd__dfxtp_2 s862 (.CLK(clknet_4_0_0_clk),
    .D(net120),
    .Q(net655));
 sky130_fd_sc_hd__dfxtp_2 s863 (.CLK(clknet_4_1_0_clk),
    .D(net126),
    .Q(net855));
 sky130_fd_sc_hd__dfxtp_1 s864 (.CLK(clknet_4_1_0_clk),
    .D(net127),
    .Q(net656));
 sky130_fd_sc_hd__dlclkp_1 s865 (.CLK(clknet_4_1_0_clk),
    .GATE(net128),
    .GCLK(net657));
 sky130_fd_sc_hd__dlclkp_2 s866 (.CLK(clknet_4_4_0_clk),
    .GATE(net143),
    .GCLK(net658));
 sky130_fd_sc_hd__dlclkp_4 s867 (.CLK(clknet_4_4_0_clk),
    .GATE(net144),
    .GCLK(net659));
 sky130_fd_sc_hd__dlxbn_1 s868 (.D(net172),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net661),
    .Q_N(net660));
 sky130_fd_sc_hd__dlxbn_2 s869 (.D(net180),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net663),
    .Q_N(net662));
 sky130_fd_sc_hd__dlxbp_1 s870 (.D(net187),
    .GATE(clknet_4_7_0_clk),
    .Q(net827),
    .Q_N(net664));
 sky130_fd_sc_hd__dlxtn_2 s871 (.D(net201),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net665));
 sky130_fd_sc_hd__dlxtn_2 s872 (.D(net207),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net666));
 sky130_fd_sc_hd__dlxtn_1 s873 (.D(net232),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net667));
 sky130_fd_sc_hd__dlxtp_1 s874 (.D(net235),
    .GATE(clknet_4_0_0_clk),
    .Q(net668));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s875 (.D(net244),
    .SLEEP_B(clknet_4_4_0_clk),
    .Q(net669));
 sky130_fd_sc_hd__dfxbp_2 s876 (.CLK(clknet_4_12_0_clk),
    .D(net281),
    .Q(net822),
    .Q_N(net670));
 sky130_fd_sc_hd__dfxbp_2 s877 (.CLK(clknet_4_9_0_clk),
    .D(net282),
    .Q(net672),
    .Q_N(net671));
 sky130_fd_sc_hd__dfxtp_1 s878 (.CLK(clknet_4_13_0_clk),
    .D(net283),
    .Q(net673));
 sky130_fd_sc_hd__dfxtp_2 s879 (.CLK(clknet_4_12_0_clk),
    .D(net289),
    .Q(net674));
 sky130_fd_sc_hd__dfxtp_1 s880 (.CLK(clknet_4_13_0_clk),
    .D(net293),
    .Q(net675));
 sky130_fd_sc_hd__dlclkp_1 s881 (.CLK(clknet_4_14_0_clk),
    .GATE(net295),
    .GCLK(net676));
 sky130_fd_sc_hd__dlclkp_2 s882 (.CLK(clknet_4_13_0_clk),
    .GATE(net297),
    .GCLK(net677));
 sky130_fd_sc_hd__dlclkp_4 s883 (.CLK(clknet_4_14_0_clk),
    .GATE(net299),
    .GCLK(net678));
 sky130_fd_sc_hd__dlxbn_1 s884 (.D(net306),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net680),
    .Q_N(net679));
 sky130_fd_sc_hd__dlxbn_1 s885 (.D(net311),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net828),
    .Q_N(net681));
 sky130_fd_sc_hd__dlxbp_1 s886 (.D(net318),
    .GATE(clknet_4_15_0_clk),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__dlxtn_1 s887 (.D(net320),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net835));
 sky130_fd_sc_hd__dlxtn_2 s888 (.D(net321),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net684));
 sky130_fd_sc_hd__dlxtn_2 s889 (.D(net322),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net850));
 sky130_fd_sc_hd__dlxtp_1 s890 (.D(net323),
    .GATE(clknet_4_15_0_clk),
    .Q(net685));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s891 (.D(net324),
    .SLEEP_B(clknet_4_15_0_clk),
    .Q(net686));
 sky130_fd_sc_hd__dfxbp_1 s892 (.CLK(clknet_4_14_0_clk),
    .D(net328),
    .Q(net818),
    .Q_N(net687));
 sky130_fd_sc_hd__dfxbp_1 s893 (.CLK(clknet_4_2_0_clk),
    .D(net344),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__dfxtp_2 s894 (.CLK(clknet_4_2_0_clk),
    .D(net346),
    .Q(net690));
 sky130_fd_sc_hd__dfxtp_2 s895 (.CLK(clknet_4_9_0_clk),
    .D(net364),
    .Q(net691));
 sky130_fd_sc_hd__dfxtp_1 s896 (.CLK(clknet_4_3_0_clk),
    .D(net367),
    .Q(net692));
 sky130_fd_sc_hd__dlclkp_1 s897 (.CLK(clknet_4_3_0_clk),
    .GATE(net370),
    .GCLK(net693));
 sky130_fd_sc_hd__dlclkp_2 s898 (.CLK(clknet_4_9_0_clk),
    .GATE(net373),
    .GCLK(net694));
 sky130_fd_sc_hd__dlclkp_4 s899 (.CLK(clknet_4_9_0_clk),
    .GATE(net393),
    .GCLK(net695));
 sky130_fd_sc_hd__dlxbn_1 s900 (.D(net398),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net697),
    .Q_N(net696));
 sky130_fd_sc_hd__dlxbn_1 s901 (.D(net403),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net816),
    .Q_N(net698));
 sky130_fd_sc_hd__dlxbp_1 s902 (.D(net406),
    .GATE(clknet_4_11_0_clk),
    .Q(net700),
    .Q_N(net699));
 sky130_fd_sc_hd__dlxtn_2 s903 (.D(net408),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net814));
 sky130_fd_sc_hd__dlxtn_1 s904 (.D(net430),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net701));
 sky130_fd_sc_hd__dlxtn_2 s905 (.D(net434),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net702));
 sky130_fd_sc_hd__dlxtp_1 s906 (.D(net493),
    .GATE(clknet_4_8_0_clk),
    .Q(net703));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s907 (.D(net499),
    .SLEEP_B(clknet_4_8_0_clk),
    .Q(net704));
 sky130_fd_sc_hd__dfxbp_1 s908 (.CLK(clknet_4_10_0_clk),
    .D(net507),
    .Q(net706),
    .Q_N(net705));
 sky130_fd_sc_hd__dfxbp_1 s909 (.CLK(clknet_4_8_0_clk),
    .D(net508),
    .Q(net708),
    .Q_N(net707));
 sky130_fd_sc_hd__dfxtp_2 s910 (.CLK(clknet_4_10_0_clk),
    .D(net511),
    .Q(net709));
 sky130_fd_sc_hd__dfxtp_1 s911 (.CLK(clknet_4_11_0_clk),
    .D(net531),
    .Q(net710));
 sky130_fd_sc_hd__dfxtp_4 s912 (.CLK(clknet_4_11_0_clk),
    .D(net532),
    .Q(net711));
 sky130_fd_sc_hd__dlclkp_1 s913 (.CLK(clknet_4_10_0_clk),
    .GATE(net545),
    .GCLK(net712));
 sky130_fd_sc_hd__dlclkp_2 s914 (.CLK(clknet_4_12_0_clk),
    .GATE(net552),
    .GCLK(net713));
 sky130_fd_sc_hd__dlclkp_4 s915 (.CLK(clknet_4_3_0_clk),
    .GATE(net558),
    .GCLK(net714));
 sky130_fd_sc_hd__dlxbn_1 s916 (.D(net562),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net716),
    .Q_N(net715));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(in0),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net718));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net719));
 sky130_fd_sc_hd__buf_1 input4 (.A(in11),
    .X(net720));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net721));
 sky130_fd_sc_hd__buf_12 input6 (.A(in13),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net723));
 sky130_fd_sc_hd__buf_4 input8 (.A(in15),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(in16),
    .X(net725));
 sky130_fd_sc_hd__buf_1 input10 (.A(in17),
    .X(net726));
 sky130_fd_sc_hd__buf_1 input11 (.A(in18),
    .X(net727));
 sky130_fd_sc_hd__buf_2 input12 (.A(in19),
    .X(net728));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(in20),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(in21),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(in22),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in23),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net734));
 sky130_fd_sc_hd__buf_1 input19 (.A(in25),
    .X(net735));
 sky130_fd_sc_hd__buf_1 input20 (.A(in26),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in28),
    .X(net738));
 sky130_fd_sc_hd__buf_2 input23 (.A(in29),
    .X(net739));
 sky130_fd_sc_hd__buf_2 input24 (.A(in3),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net741));
 sky130_fd_sc_hd__buf_2 input26 (.A(in31),
    .X(net742));
 sky130_fd_sc_hd__buf_4 input27 (.A(in32),
    .X(net743));
 sky130_fd_sc_hd__buf_4 input28 (.A(in33),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(in34),
    .X(net745));
 sky130_fd_sc_hd__buf_1 input30 (.A(in35),
    .X(net746));
 sky130_fd_sc_hd__buf_2 input31 (.A(in36),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(in37),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_8 input33 (.A(in38),
    .X(net749));
 sky130_fd_sc_hd__buf_1 input34 (.A(in39),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(in4),
    .X(net751));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net752));
 sky130_fd_sc_hd__buf_2 input37 (.A(in41),
    .X(net753));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net754));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(in43),
    .X(net755));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net756));
 sky130_fd_sc_hd__buf_1 input41 (.A(in46),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(in47),
    .X(net758));
 sky130_fd_sc_hd__buf_1 input43 (.A(in48),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in49),
    .X(net760));
 sky130_fd_sc_hd__buf_1 input45 (.A(in5),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(in50),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(in51),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(in52),
    .X(net764));
 sky130_fd_sc_hd__buf_1 input49 (.A(in53),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in54),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(in57),
    .X(net767));
 sky130_fd_sc_hd__buf_1 input52 (.A(in58),
    .X(net768));
 sky130_fd_sc_hd__buf_1 input53 (.A(in59),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_8 input54 (.A(in6),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(in60),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(in61),
    .X(net772));
 sky130_fd_sc_hd__buf_1 input57 (.A(in62),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(in63),
    .X(net774));
 sky130_fd_sc_hd__buf_1 input59 (.A(in64),
    .X(net775));
 sky130_fd_sc_hd__buf_1 input60 (.A(in65),
    .X(net776));
 sky130_fd_sc_hd__buf_1 input61 (.A(in66),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(in67),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_4 input63 (.A(in68),
    .X(net779));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(in69),
    .X(net780));
 sky130_fd_sc_hd__buf_1 input65 (.A(in7),
    .X(net781));
 sky130_fd_sc_hd__buf_2 input66 (.A(in70),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(in71),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_4 input68 (.A(in72),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(in73),
    .X(net785));
 sky130_fd_sc_hd__buf_1 input70 (.A(in74),
    .X(net786));
 sky130_fd_sc_hd__buf_1 input71 (.A(in75),
    .X(net787));
 sky130_fd_sc_hd__dlymetal6s2s_1 input72 (.A(in76),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(in77),
    .X(net789));
 sky130_fd_sc_hd__buf_1 input74 (.A(in78),
    .X(net790));
 sky130_fd_sc_hd__buf_2 input75 (.A(in79),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(in8),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(in80),
    .X(net793));
 sky130_fd_sc_hd__buf_1 input78 (.A(in81),
    .X(net794));
 sky130_fd_sc_hd__buf_1 input79 (.A(in82),
    .X(net795));
 sky130_fd_sc_hd__buf_1 input80 (.A(in83),
    .X(net796));
 sky130_fd_sc_hd__buf_1 input81 (.A(in84),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(in85),
    .X(net798));
 sky130_fd_sc_hd__buf_1 input83 (.A(in86),
    .X(net799));
 sky130_fd_sc_hd__buf_4 input84 (.A(in87),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(in88),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(in89),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(in9),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_4 input88 (.A(in90),
    .X(net804));
 sky130_fd_sc_hd__buf_1 input89 (.A(in91),
    .X(net805));
 sky130_fd_sc_hd__buf_2 input90 (.A(in92),
    .X(net806));
 sky130_fd_sc_hd__buf_1 input91 (.A(in93),
    .X(net807));
 sky130_fd_sc_hd__buf_1 input92 (.A(in94),
    .X(net808));
 sky130_fd_sc_hd__buf_1 input93 (.A(in95),
    .X(net809));
 sky130_fd_sc_hd__buf_1 input94 (.A(in96),
    .X(net810));
 sky130_fd_sc_hd__buf_4 input95 (.A(in97),
    .X(net811));
 sky130_fd_sc_hd__buf_1 input96 (.A(in98),
    .X(net812));
 sky130_fd_sc_hd__dlymetal6s2s_1 input97 (.A(in99),
    .X(net813));
 sky130_fd_sc_hd__buf_2 output98 (.A(net814),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(clknet_1_1__leaf_net815),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output100 (.A(net816),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output101 (.A(net817),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output102 (.A(net818),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output103 (.A(net819),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net820),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(clknet_1_1__leaf_net821),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output106 (.A(net822),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net823),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net824),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output109 (.A(net825),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output110 (.A(net826),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net827),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net828),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net829),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net830),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net831),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(clknet_1_1__leaf_net832),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net833),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net834),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net835),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_4 output120 (.A(net836),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net837),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_4 output122 (.A(net954),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output123 (.A(net839),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output124 (.A(net840),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net841),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net842),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net843),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(clknet_1_1__leaf_net844),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net845),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_4 output130 (.A(net846),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net847),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_4 output132 (.A(net848),
    .X(out48));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net849),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output134 (.A(net850),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_4 output135 (.A(net851),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output136 (.A(net852),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_4 output137 (.A(net853),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output138 (.A(net854),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output139 (.A(net855),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net898),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net857),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(clknet_1_1__leaf_net858),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net859),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_4 output144 (.A(net860),
    .X(out61));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net861),
    .X(out62));
 sky130_fd_sc_hd__clkbuf_4 output146 (.A(net934),
    .X(out65));
 sky130_fd_sc_hd__buf_2 output147 (.A(net863),
    .X(out68));
 sky130_fd_sc_hd__buf_2 output148 (.A(net864),
    .X(out69));
 sky130_fd_sc_hd__buf_2 output149 (.A(net865),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net866),
    .X(out73));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net867),
    .X(out76));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net868),
    .X(out79));
 sky130_fd_sc_hd__buf_2 output153 (.A(net869),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net870),
    .X(out82));
 sky130_fd_sc_hd__clkbuf_4 output155 (.A(net871),
    .X(out83));
 sky130_fd_sc_hd__buf_2 output156 (.A(net872),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output157 (.A(net873),
    .X(out87));
 sky130_fd_sc_hd__clkbuf_4 output158 (.A(net874),
    .X(out89));
 sky130_fd_sc_hd__buf_2 output159 (.A(net875),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 output160 (.A(net876),
    .X(out91));
 sky130_fd_sc_hd__clkbuf_4 output161 (.A(net877),
    .X(out92));
 sky130_fd_sc_hd__clkbuf_4 output162 (.A(net878),
    .X(out93));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net879),
    .X(out94));
 sky130_fd_sc_hd__clkbuf_4 output164 (.A(net880),
    .X(out96));
 sky130_fd_sc_hd__clkbuf_4 output165 (.A(net881),
    .X(out97));
 sky130_fd_sc_hd__buf_1 wire166 (.A(net976),
    .X(net882));
 sky130_fd_sc_hd__buf_1 max_cap167 (.A(net884),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_2 wire168 (.A(net977),
    .X(net884));
 sky130_fd_sc_hd__buf_2 fanout169 (.A(net886),
    .X(net885));
 sky130_fd_sc_hd__buf_2 fanout170 (.A(net887),
    .X(net886));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net110),
    .X(net887));
 sky130_fd_sc_hd__buf_2 wire172 (.A(net55),
    .X(net888));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net891),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_4 fanout174 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_2 fanout175 (.A(net335),
    .X(net891));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(net142),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_4 fanout178 (.A(net142),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_4 fanout179 (.A(net107),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_2 max_cap180 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_2 max_cap181 (.A(net978),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_2 max_cap182 (.A(net899),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_2 max_cap183 (.A(net856),
    .X(net899));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap184 (.A(net901),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_2 max_cap185 (.A(net860),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_1 max_cap186 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__buf_1 max_cap187 (.A(net979),
    .X(net903));
 sky130_fd_sc_hd__buf_1 max_cap188 (.A(net980),
    .X(net904));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net449),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_1 max_cap190 (.A(net492),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_2 max_cap191 (.A(net278),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net153),
    .X(net908));
 sky130_fd_sc_hd__buf_12 fanout193 (.A(net11),
    .X(net909));
 sky130_fd_sc_hd__clkbuf_2 max_cap194 (.A(net268),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_2 max_cap195 (.A(net51),
    .X(net911));
 sky130_fd_sc_hd__clkbuf_2 max_cap196 (.A(net38),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_2 max_cap197 (.A(net874),
    .X(net913));
 sky130_fd_sc_hd__buf_4 fanout198 (.A(net377),
    .X(net914));
 sky130_fd_sc_hd__buf_2 fanout199 (.A(net331),
    .X(net915));
 sky130_fd_sc_hd__buf_1 max_cap200 (.A(net174),
    .X(net916));
 sky130_fd_sc_hd__clkbuf_2 max_cap201 (.A(net52),
    .X(net917));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net28),
    .X(net918));
 sky130_fd_sc_hd__buf_1 max_cap203 (.A(net1),
    .X(net919));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(net701),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_8 fanout205 (.A(net691),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_4 wire206 (.A(net668),
    .X(net922));
 sky130_fd_sc_hd__buf_4 max_cap207 (.A(net166),
    .X(net923));
 sky130_fd_sc_hd__buf_4 fanout208 (.A(net47),
    .X(net924));
 sky130_fd_sc_hd__buf_2 fanout209 (.A(net47),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_8 fanout210 (.A(net6),
    .X(net926));
 sky130_fd_sc_hd__buf_12 fanout211 (.A(net722),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_8 fanout212 (.A(net718),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_8 fanout213 (.A(net729),
    .X(net929));
 sky130_fd_sc_hd__clkinv_1 c534_1 (.A(clknet_1_1__leaf_net714),
    .Y(net930));
 sky130_fd_sc_hd__clkinv_1 net899_2 (.A(clknet_1_0__leaf_net714),
    .Y(net931));
 sky130_fd_sc_hd__clkinv_1 net899_3 (.A(clknet_1_1__leaf_net714),
    .Y(net932));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net714 (.A(net714),
    .X(clknet_0_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net714 (.A(clknet_0_net714),
    .X(clknet_1_0__leaf_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net714 (.A(clknet_0_net714),
    .X(clknet_1_1__leaf_net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net360 (.A(net360),
    .X(clknet_0_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net360 (.A(clknet_0_net360),
    .X(clknet_1_0__leaf_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net360 (.A(clknet_0_net360),
    .X(clknet_1_1__leaf_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net410 (.A(net410),
    .X(clknet_0_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_0__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_1__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net404 (.A(net404),
    .X(clknet_0_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net378 (.A(net378),
    .X(clknet_0_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_1__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net417 (.A(net417),
    .X(clknet_0_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net417 (.A(clknet_0_net417),
    .X(clknet_1_0__leaf_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net417 (.A(clknet_0_net417),
    .X(clknet_1_1__leaf_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net627 (.A(net627),
    .X(clknet_0_net627));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net627 (.A(clknet_0_net627),
    .X(clknet_1_0__leaf_net627));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net627 (.A(clknet_0_net627),
    .X(clknet_1_1__leaf_net627));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net333 (.A(net333),
    .X(clknet_0_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net333 (.A(clknet_0_net333),
    .X(clknet_1_0__leaf_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net333 (.A(clknet_0_net333),
    .X(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net355 (.A(net355),
    .X(clknet_0_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net355 (.A(net956),
    .X(clknet_1_0__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_1__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net477 (.A(net477),
    .X(clknet_0_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net477 (.A(clknet_0_net477),
    .X(clknet_1_0__leaf_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net477 (.A(clknet_0_net477),
    .X(clknet_1_1__leaf_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net361 (.A(net361),
    .X(clknet_0_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net368 (.A(net368),
    .X(clknet_0_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_0__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_1__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net694 (.A(net694),
    .X(clknet_0_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net381 (.A(net381),
    .X(clknet_0_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_0__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_1__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net858 (.A(net858),
    .X(clknet_0_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net858 (.A(clknet_0_net858),
    .X(clknet_1_0__leaf_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net858 (.A(clknet_0_net858),
    .X(clknet_1_1__leaf_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net371 (.A(net371),
    .X(clknet_0_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_0__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_1__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net369 (.A(net369),
    .X(clknet_0_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_0__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_1__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net359 (.A(net359),
    .X(clknet_0_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net359 (.A(clknet_0_net359),
    .X(clknet_1_0__leaf_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net359 (.A(clknet_0_net359),
    .X(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net382 (.A(net382),
    .X(clknet_0_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_0__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_1__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net383 (.A(net383),
    .X(clknet_0_net383));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net383 (.A(clknet_0_net383),
    .X(clknet_1_0__leaf_net383));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net383 (.A(clknet_0_net383),
    .X(clknet_1_1__leaf_net383));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net695 (.A(net695),
    .X(clknet_0_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net695 (.A(clknet_0_net695),
    .X(clknet_1_0__leaf_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net695 (.A(clknet_0_net695),
    .X(clknet_1_1__leaf_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net395 (.A(net395),
    .X(clknet_0_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net395 (.A(clknet_0_net395),
    .X(clknet_1_0__leaf_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net395 (.A(clknet_0_net395),
    .X(clknet_1_1__leaf_net395));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net832 (.A(net832),
    .X(clknet_0_net832));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net832 (.A(clknet_0_net832),
    .X(clknet_1_0__leaf_net832));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net832 (.A(clknet_0_net832),
    .X(clknet_1_1__leaf_net832));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net815 (.A(net815),
    .X(clknet_0_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net815 (.A(clknet_0_net815),
    .X(clknet_1_0__leaf_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net815 (.A(clknet_0_net815),
    .X(clknet_1_1__leaf_net815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net435 (.A(net435),
    .X(clknet_0_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_0__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net693 (.A(net693),
    .X(clknet_0_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net484 (.A(net484),
    .X(clknet_0_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net484 (.A(clknet_0_net484),
    .X(clknet_1_0__leaf_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net484 (.A(clknet_0_net484),
    .X(clknet_1_1__leaf_net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net365 (.A(net365),
    .X(clknet_0_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net713 (.A(net713),
    .X(clknet_0_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net713 (.A(clknet_0_net713),
    .X(clknet_1_0__leaf_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net713 (.A(clknet_0_net713),
    .X(clknet_1_1__leaf_net713));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net821 (.A(net821),
    .X(clknet_0_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net821 (.A(clknet_0_net821),
    .X(clknet_1_0__leaf_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net821 (.A(clknet_0_net821),
    .X(clknet_1_1__leaf_net821));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net712 (.A(net712),
    .X(clknet_0_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_0__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net712 (.A(clknet_0_net712),
    .X(clknet_1_1__leaf_net712));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net678 (.A(net678),
    .X(clknet_0_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net678 (.A(clknet_0_net678),
    .X(clknet_1_0__leaf_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net678 (.A(clknet_0_net678),
    .X(clknet_1_1__leaf_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net305 (.A(net305),
    .X(clknet_0_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_0__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_1__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net677 (.A(net677),
    .X(clknet_0_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_0__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net677 (.A(clknet_0_net677),
    .X(clknet_1_1__leaf_net677));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net676 (.A(net676),
    .X(clknet_0_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_0__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_1__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net302 (.A(net302),
    .X(clknet_0_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_0__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_1__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net307 (.A(net307),
    .X(clknet_0_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_0__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_1__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net296 (.A(net296),
    .X(clknet_0_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_0__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_1__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net298 (.A(net298),
    .X(clknet_0_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_0__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_1__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net659 (.A(net659),
    .X(clknet_0_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net659 (.A(clknet_0_net659),
    .X(clknet_1_0__leaf_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net659 (.A(clknet_0_net659),
    .X(clknet_1_1__leaf_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net202 (.A(net202),
    .X(clknet_0_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_0__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net202 (.A(clknet_0_net202),
    .X(clknet_1_1__leaf_net202));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net182 (.A(net182),
    .X(clknet_0_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net425 (.A(net425),
    .X(clknet_0_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_0__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_1__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net424 (.A(net424),
    .X(clknet_0_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net424 (.A(clknet_0_net424),
    .X(clknet_1_0__leaf_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net424 (.A(clknet_0_net424),
    .X(clknet_1_1__leaf_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net314 (.A(net314),
    .X(clknet_0_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net314 (.A(clknet_0_net314),
    .X(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net314 (.A(clknet_0_net314),
    .X(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net317 (.A(net317),
    .X(clknet_0_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_0__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_1__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net287 (.A(net287),
    .X(clknet_0_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_0__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_1__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net294 (.A(net294),
    .X(clknet_0_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net206 (.A(net206),
    .X(clknet_0_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net206 (.A(clknet_0_net206),
    .X(clknet_1_0__leaf_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net206 (.A(clknet_0_net206),
    .X(clknet_1_1__leaf_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net195 (.A(net195),
    .X(clknet_0_net195));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net195 (.A(clknet_0_net195),
    .X(clknet_1_0__leaf_net195));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net195 (.A(clknet_0_net195),
    .X(clknet_1_1__leaf_net195));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net316 (.A(net316),
    .X(clknet_0_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_0__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_1__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net192 (.A(net192),
    .X(clknet_0_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net192 (.A(clknet_0_net192),
    .X(clknet_1_0__leaf_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net192 (.A(clknet_0_net192),
    .X(clknet_1_1__leaf_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net844 (.A(net844),
    .X(clknet_0_net844));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net844 (.A(clknet_0_net844),
    .X(clknet_1_0__leaf_net844));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net844 (.A(clknet_0_net844),
    .X(clknet_1_1__leaf_net844));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net184 (.A(net184),
    .X(clknet_0_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net184 (.A(clknet_0_net184),
    .X(clknet_1_0__leaf_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net184 (.A(clknet_0_net184),
    .X(clknet_1_1__leaf_net184));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net288 (.A(net288),
    .X(clknet_0_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_1__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net285 (.A(net285),
    .X(clknet_0_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_0__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_1__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net286 (.A(net286),
    .X(clknet_0_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_0__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_1__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net183 (.A(net183),
    .X(clknet_0_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_0__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net183 (.A(clknet_0_net183),
    .X(clknet_1_1__leaf_net183));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net165 (.A(net165),
    .X(clknet_0_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net167 (.A(net167),
    .X(clknet_0_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_0__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_1__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net625 (.A(net625),
    .X(clknet_0_net625));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net625 (.A(clknet_0_net625),
    .X(clknet_1_0__leaf_net625));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net625 (.A(clknet_0_net625),
    .X(clknet_1_1__leaf_net625));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net151 (.A(net151),
    .X(clknet_0_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net151 (.A(clknet_0_net151),
    .X(clknet_1_0__leaf_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net151 (.A(clknet_0_net151),
    .X(clknet_1_1__leaf_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net150 (.A(net150),
    .X(clknet_0_net150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net150 (.A(clknet_0_net150),
    .X(clknet_1_0__leaf_net150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net150 (.A(clknet_0_net150),
    .X(clknet_1_1__leaf_net150));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net156 (.A(net156),
    .X(clknet_0_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net154 (.A(net154),
    .X(clknet_0_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net154 (.A(clknet_0_net154),
    .X(clknet_1_0__leaf_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net154 (.A(clknet_0_net154),
    .X(clknet_1_1__leaf_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net161 (.A(net161),
    .X(clknet_0_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net159 (.A(net159),
    .X(clknet_0_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_0__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_1__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net157 (.A(net157),
    .X(clknet_0_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_1__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net658 (.A(net658),
    .X(clknet_0_net658));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net658 (.A(clknet_0_net658),
    .X(clknet_1_0__leaf_net658));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net658 (.A(clknet_0_net658),
    .X(clknet_1_1__leaf_net658));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net245 (.A(net245),
    .X(clknet_0_net245));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net245 (.A(clknet_0_net245),
    .X(clknet_1_0__leaf_net245));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net245 (.A(clknet_0_net245),
    .X(clknet_1_1__leaf_net245));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net657 (.A(net657),
    .X(clknet_0_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_0__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_1__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net219 (.A(net219),
    .X(clknet_0_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net231 (.A(net231),
    .X(clknet_0_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net231 (.A(clknet_0_net231),
    .X(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net231 (.A(clknet_0_net231),
    .X(clknet_1_1__leaf_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net223 (.A(net223),
    .X(clknet_0_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_0__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_1__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net229 (.A(net229),
    .X(clknet_0_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net229 (.A(clknet_0_net229),
    .X(clknet_1_0__leaf_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net229 (.A(clknet_0_net229),
    .X(clknet_1_1__leaf_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net228 (.A(net228),
    .X(clknet_0_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_0__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_1__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net220 (.A(net220),
    .X(clknet_0_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net337 (.A(net337),
    .X(clknet_0_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net337 (.A(clknet_0_net337),
    .X(clknet_1_0__leaf_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net337 (.A(clknet_0_net337),
    .X(clknet_1_1__leaf_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net212 (.A(net212),
    .X(clknet_0_net212));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net212 (.A(clknet_0_net212),
    .X(clknet_1_0__leaf_net212));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net212 (.A(clknet_0_net212),
    .X(clknet_1_1__leaf_net212));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net862),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net336),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net933),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net862),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net935),
    .X(net936));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer6 (.A(net936),
    .X(net937));
 sky130_fd_sc_hd__buf_4 rebuffer7 (.A(net18),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net938),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net17),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net20),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net941),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net11),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net358),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net944),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net944),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net946),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net944),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net24),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net949),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net949),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net24),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net24),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net838),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net81),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(clknet_0_net355),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net218),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net957),
    .X(net958));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer28 (.A(net958),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(clknet_1_1__leaf_net359),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net586),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net459),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net269),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net846),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net703),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net353),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net600),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net665),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net668),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net630),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net690),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net692),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net647),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net270),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net214),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_1 wire1 (.A(net194),
    .X(net976));
 sky130_fd_sc_hd__buf_1 wire2 (.A(net138),
    .X(net977));
 sky130_fd_sc_hd__buf_1 max_cap3 (.A(net48),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_1 wire4 (.A(net496),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_1 wire5 (.A(net4),
    .X(net980));
 sky130_fd_sc_hd__buf_6 max_cap6 (.A(net7),
    .X(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_C (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_C (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_D (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_Y (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A3 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_C (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_D1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_RESET_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_Q_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_Q (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_D (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_Q (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_D (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_Q (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_Q_N (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_C (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A_N (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_Q (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_RESET_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_Y (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_S1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A_N (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A3 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_C_N (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_X (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B_N (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_Y (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_C1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_Q_N (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_C_N (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_Q (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_Y (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net156_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A_N (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A0 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_X (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A0 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A0 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_SCD (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_X (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A0 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A_N (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_Y (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_C (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_C1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer26_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_C (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_S0 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S0 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SCE (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_Q_N (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_RESET_B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_Q (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A_N (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_C (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_C_N (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net231_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_Y (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_SCE (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_Y (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_C (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer21_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_C (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_C (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCE (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_Q (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A3 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A_N (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_SCE (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_D (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_Q_N (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_Q (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_C (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCD (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_C (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_C1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_X (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_C1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_D (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S0 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_C (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_X (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_Q (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_Y (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A0 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_Q (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_D1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_Q_N (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_Q (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_C (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_Y (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SCE (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_Y (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_SCE (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_Q (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A3 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_Y (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_C1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_Y (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_C1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_X (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_RESET_B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_SCD (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_S0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_DE (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_Y (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_B1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_D1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_Q_N (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_Q (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_Q (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_B1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A0 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A3 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_X (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_Y (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_SCE (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_D (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_D (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SCD (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_D (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_SCD (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A2 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_X (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_C1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_C1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_Q_N (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A0 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_B1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_C (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_Q (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap195_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_Y (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_C1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_Q_N (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_X (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_D (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_D (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_Y (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_Q (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_S1 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S1 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_SCE (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_SCE (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_SET_B (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_Q (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_D1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_SCE (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_Q (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_S1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_D1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S0 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_C1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_D1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_C (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_C (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_C (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_C (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_D_N (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_C (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_D1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_Q (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_C (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_C1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_Q (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_S1 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_C1 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_D (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_D (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_Q (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_Q (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_D1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_Q (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SCE (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_D1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_Q (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_Q_N (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A3 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_Q_N (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_C (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_D (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_Q (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_C1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S0 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_Q (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_S1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_B (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_SET_B (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_Q_N (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_D1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_Q (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_D1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_D (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_Q (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_D1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_D1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold38_A (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire206_A (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_Q (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_C1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_D1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_Q_N (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_S1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_C (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_Q_N (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SET_B (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_D1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_D (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_Q (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_D1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_C (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_Q (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_D1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_C (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_D1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_C1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_s895_Q (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_Y (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_Q (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_SCE (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A3 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_D (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_C1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_C1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_D1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_SCD (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_C1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_C1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A3 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_C (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_D (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_C1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_B1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_D (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_D1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A_N (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_D1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_D1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_C1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_C (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B_N (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A_N (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_C (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_S0 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_C_N (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_C1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B_N (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A0 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_C_N (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_C (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_RESET_B (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_C (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_C (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A0 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_C_N (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_C (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SCD (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_C1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A3 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A0 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_B1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_C (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_C1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_X (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_RESET_B (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_D1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_C (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_C1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A2 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_X (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_S0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A2 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_B1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_B1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_B (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_X (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_C1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_B (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_C1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_D1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_D1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_C1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S0 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_C1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_C1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_B1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_Q (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_D1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_Q (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_Q (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_D1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_B1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_Q (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_C1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_B1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_SCE (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_Q (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_Q (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_D1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_D (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_Y (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net832_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_D1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_D1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_Q_N (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_SCE (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold33_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_Q (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_C_N (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_Q (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_C1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_D (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_Q (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_B1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_D (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_Y (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_Q (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_C1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_S0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_Y (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_X (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A3 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B_N (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_Q (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_D1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_Y (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_RESET_B (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_D1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_D_N (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap197_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_Y (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_Q (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_S1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_C1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_X (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_B1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SET_B (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire172_X (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_D1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_D_N (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_D1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_D (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_B1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_SCD (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_D_N (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_C1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_SCE (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_SET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_B1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_D1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_C (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_C (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_C1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_C1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_SCE (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_C_N (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCE (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_C (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_C1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_D (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_D1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C_N (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_C_N (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_C1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_C (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_C (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_SCD (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_C_N (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_C (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap180_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap181_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap180_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap182_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_C (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_SCD (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_SCD (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_C1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCE (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_C (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_RESET_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_SET_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_C_N (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap194_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A2 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_C1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_C1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_D1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_C (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_C (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_C1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_B1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_S0 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_C_N (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_D_N (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A_N (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_C (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_D1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_C1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_SET_B (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire206_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_D1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCE (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap207_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_C (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_S0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_C (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_C_N (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_D1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_C1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_RESET_B (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_D1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_D1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_C1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_B (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_B1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_C_N (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_C_N (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_C (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_C1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_SCD (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_C (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_C (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_C (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_SLEEP_B (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_B1 (.DIODE(clknet_1_1__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_S1 (.DIODE(clknet_1_1__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(clknet_1_1__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net832_X (.DIODE(clknet_1_1__leaf_net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_C (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S1 (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_C1 (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S1 (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_C (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B1 (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B1 (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_D1 (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_D1 (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net182_X (.DIODE(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_C (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCD (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_SCE (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net182_X (.DIODE(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(clknet_1_1__leaf_net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_D (.DIODE(clknet_1_1__leaf_net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(clknet_1_1__leaf_net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(clknet_1_1__leaf_net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net844_X (.DIODE(clknet_1_1__leaf_net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(clknet_1_1__leaf_net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S1 (.DIODE(clknet_1_1__leaf_net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(clknet_1_1__leaf_net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net625_X (.DIODE(clknet_1_1__leaf_net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net156_A (.DIODE(clknet_0_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net156_A (.DIODE(clknet_0_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net156_X (.DIODE(clknet_0_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_S0 (.DIODE(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_S1 (.DIODE(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net156_X (.DIODE(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCD (.DIODE(clknet_1_0__leaf_net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A1 (.DIODE(clknet_1_0__leaf_net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_SCD (.DIODE(clknet_1_0__leaf_net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_SCE (.DIODE(clknet_1_0__leaf_net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A1 (.DIODE(clknet_1_0__leaf_net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A2 (.DIODE(clknet_1_0__leaf_net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net245_X (.DIODE(clknet_1_0__leaf_net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net231_A (.DIODE(clknet_0_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net231_A (.DIODE(clknet_0_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net231_X (.DIODE(clknet_0_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SET_B (.DIODE(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S1 (.DIODE(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A1 (.DIODE(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A1 (.DIODE(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net231_X (.DIODE(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_SET_B (.DIODE(clknet_1_1__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(clknet_1_1__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A1 (.DIODE(clknet_1_1__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_B1 (.DIODE(clknet_1_1__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net231_X (.DIODE(clknet_1_1__leaf_net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_B1 (.DIODE(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A3 (.DIODE(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A0 (.DIODE(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net220_X (.DIODE(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_B1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_C_N (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net929));
 sky130_fd_sc_hd__or4bb_1 clone1 (.A(net751),
    .B(net981),
    .C_N(net991),
    .D_N(net8),
    .X(net982));
 sky130_fd_sc_hd__a2111o_1 clone2 (.A1(net20),
    .A2(net10),
    .B1(net981),
    .C1(net984),
    .D1(net12),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net21),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer31 (.A(net23),
    .X(net985));
 sky130_fd_sc_hd__buf_8 rebuffer32 (.A(net23),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net986),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_1 clone34 (.A(net722),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_1 clone35 (.A(net11),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_1 clone36 (.A(net11),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_1 clone37 (.A(net722),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer38 (.A(net722),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net992),
    .X(net993));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
endmodule
